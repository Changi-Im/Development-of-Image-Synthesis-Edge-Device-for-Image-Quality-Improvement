module database_pixel(clk,datata,re,address,we,dp,address_p);

	parameter SIZE=0;

	input 							clk; 		// clock
	output	reg	signed	[SIZE-1:0]	datata;		// read data
	input 							re,we; 		// read signal, write signal 
	input 				[15:0] 		address;	// read address from database_pixel to RAM
	input 		signed 	[SIZE-1:0] 	dp; 		// write data from testbench to database_pixel
	input 				[15:0] 		address_p;	// write address


   
	reg signed [SIZE-1:0] storage [0:3199];

	initial begin
storage[0] = 0;
storage[1] = 0;
storage[2] = 0;
storage[3] = 0;
storage[4] = 0;
storage[5] = 0;
storage[6] = 0;
storage[7] = 0;
storage[8] = 0;
storage[9] = 0;
storage[10] = 0;
storage[11] = 0;
storage[12] = 0;
storage[13] = 0;
storage[14] = 0;
storage[15] = 0;
storage[16] = 0;
storage[17] = 0;
storage[18] = 0;
storage[19] = 0;
storage[20] = 0;
storage[21] = 0;
storage[22] = 0;
storage[23] = 0;
storage[24] = 0;
storage[25] = 0;
storage[26] = 0;
storage[27] = 0;
storage[28] = 0;
storage[29] = 0;
storage[30] = 0;
storage[31] = 0;
storage[32] = 0;
storage[33] = 0;
storage[34] = 0;
storage[35] = 0;
storage[36] = 0;
storage[37] = 0;
storage[38] = 0;
storage[39] = 0;
storage[40] = 0;
storage[41] = 0;
storage[42] = 0;
storage[43] = 0;
storage[44] = 0;
storage[45] = 0;
storage[46] = 0;
storage[47] = 0;
storage[48] = 0;
storage[49] = 0;
storage[50] = 0;
storage[51] = 0;
storage[52] = 0;
storage[53] = 0;
storage[54] = 0;
storage[55] = 0;
storage[56] = 0;
storage[57] = 0;
storage[58] = 0;
storage[59] = 0;
storage[60] = 0;
storage[61] = 0;
storage[62] = 0;
storage[63] = 0;
storage[64] = 0;
storage[65] = 0;
storage[66] = 0;
storage[67] = 0;
storage[68] = 0;
storage[69] = 0;
storage[70] = 0;
storage[71] = 0;
storage[72] = 0;
storage[73] = 0;
storage[74] = 0;
storage[75] = 0;
storage[76] = 0;
storage[77] = 0;
storage[78] = 0;
storage[79] = 0;
storage[80] = 0;
storage[81] = 0;
storage[82] = 0;
storage[83] = 0;
storage[84] = 0;
storage[85] = 0;
storage[86] = 0;
storage[87] = 0;
storage[88] = 0;
storage[89] = 0;
storage[90] = 0;
storage[91] = 0;
storage[92] = 0;
storage[93] = 0;
storage[94] = 0;
storage[95] = 0;
storage[96] = 0;
storage[97] = 0;
storage[98] = 0;
storage[99] = 0;
storage[100] = 0;
storage[101] = 0;
storage[102] = 0;
storage[103] = 0;
storage[104] = 0;
storage[105] = 0;
storage[106] = 0;
storage[107] = 0;
storage[108] = 0;
storage[109] = 0;
storage[110] = 0;
storage[111] = 0;
storage[112] = 0;
storage[113] = 0;
storage[114] = 0;
storage[115] = 0;
storage[116] = 0;
storage[117] = 0;
storage[118] = 0;
storage[119] = 0;
storage[120] = 0;
storage[121] = 0;
storage[122] = 0;
storage[123] = 0;
storage[124] = 0;
storage[125] = 0;
storage[126] = 0;
storage[127] = 0;
storage[128] = 0;
storage[129] = 0;
storage[130] = 0;
storage[131] = 0;
storage[132] = 0;
storage[133] = 0;
storage[134] = 0;
storage[135] = 0;
storage[136] = 0;
storage[137] = 0;
storage[138] = 0;
storage[139] = 0;
storage[140] = 0;
storage[141] = 0;
storage[142] = 0;
storage[143] = 0;
storage[144] = 0;
storage[145] = 0;
storage[146] = 0;
storage[147] = 0;
storage[148] = 0;
storage[149] = 0;
storage[150] = 0;
storage[151] = 0;
storage[152] = 0;
storage[153] = 0;
storage[154] = 0;
storage[155] = 0;
storage[156] = 0;
storage[157] = 0;
storage[158] = 0;
storage[159] = 0;
storage[160] = 0;
storage[161] = 0;
storage[162] = 0;
storage[163] = 0;
storage[164] = 0;
storage[165] = 0;
storage[166] = 0;
storage[167] = 0;
storage[168] = 0;
storage[169] = 0;
storage[170] = 0;
storage[171] = 0;
storage[172] = 0;
storage[173] = 0;
storage[174] = 0;
storage[175] = 0;
storage[176] = 0;
storage[177] = 0;
storage[178] = 0;
storage[179] = 0;
storage[180] = 0;
storage[181] = 0;
storage[182] = 0;
storage[183] = 0;
storage[184] = 0;
storage[185] = 0;
storage[186] = 0;
storage[187] = 0;
storage[188] = 0;
storage[189] = 0;
storage[190] = 0;
storage[191] = 0;
storage[192] = 0;
storage[193] = 0;
storage[194] = 0;
storage[195] = 0;
storage[196] = 0;
storage[197] = 0;
storage[198] = 0;
storage[199] = 0;
storage[200] = 0;
storage[201] = 0;
storage[202] = 0;
storage[203] = 0;
storage[204] = 0;
storage[205] = 0;
storage[206] = 0;
storage[207] = 0;
storage[208] = 0;
storage[209] = 0;
storage[210] = 0;
storage[211] = 0;
storage[212] = 0;
storage[213] = 0;
storage[214] = 0;
storage[215] = 0;
storage[216] = 0;
storage[217] = 0;
storage[218] = 0;
storage[219] = 0;
storage[220] = 0;
storage[221] = 0;
storage[222] = 0;
storage[223] = 0;
storage[224] = 0;
storage[225] = 0;
storage[226] = 0;
storage[227] = 0;
storage[228] = 0;
storage[229] = 0;
storage[230] = 0;
storage[231] = 0;
storage[232] = 0;
storage[233] = 0;
storage[234] = 0;
storage[235] = 0;
storage[236] = 0;
storage[237] = 0;
storage[238] = 0;
storage[239] = 0;
storage[240] = 0;
storage[241] = 0;
storage[242] = 0;
storage[243] = 0;
storage[244] = 0;
storage[245] = 0;
storage[246] = 0;
storage[247] = 0;
storage[248] = 0;
storage[249] = 0;
storage[250] = 0;
storage[251] = 0;
storage[252] = 0;
storage[253] = 0;
storage[254] = 0;
storage[255] = 0;
storage[256] = 0;
storage[257] = 0;
storage[258] = 0;
storage[259] = 0;
storage[260] = 0;
storage[261] = 0;
storage[262] = 0;
storage[263] = 0;
storage[264] = 0;
storage[265] = 0;
storage[266] = 0;
storage[267] = 0;
storage[268] = 0;
storage[269] = 0;
storage[270] = 0;
storage[271] = 0;
storage[272] = 0;
storage[273] = 0;
storage[274] = 0;
storage[275] = 0;
storage[276] = 0;
storage[277] = 0;
storage[278] = 0;
storage[279] = 0;
storage[280] = 0;
storage[281] = 0;
storage[282] = 0;
storage[283] = 0;
storage[284] = 0;
storage[285] = 0;
storage[286] = 0;
storage[287] = 0;
storage[288] = 0;
storage[289] = 0;
storage[290] = 0;
storage[291] = 0;
storage[292] = 0;
storage[293] = 0;
storage[294] = 0;
storage[295] = 0;
storage[296] = 0;
storage[297] = 0;
storage[298] = 0;
storage[299] = 0;
storage[300] = 0;
storage[301] = 0;
storage[302] = 0;
storage[303] = 0;
storage[304] = 0;
storage[305] = 0;
storage[306] = 0;
storage[307] = 0;
storage[308] = 0;
storage[309] = 0;
storage[310] = 0;
storage[311] = 0;
storage[312] = 0;
storage[313] = 0;
storage[314] = 0;
storage[315] = 0;
storage[316] = 0;
storage[317] = 0;
storage[318] = 0;
storage[319] = 0;
storage[320] = 0;
storage[321] = 0;
storage[322] = 0;
storage[323] = 0;
storage[324] = 0;
storage[325] = 0;
storage[326] = 0;
storage[327] = 0;
storage[328] = 0;
storage[329] = 0;
storage[330] = 0;
storage[331] = 0;
storage[332] = 0;
storage[333] = 0;
storage[334] = 0;
storage[335] = 0;
storage[336] = 0;
storage[337] = 0;
storage[338] = 0;
storage[339] = 0;
storage[340] = 0;
storage[341] = 0;
storage[342] = 0;
storage[343] = 0;
storage[344] = 0;
storage[345] = 0;
storage[346] = 0;
storage[347] = 0;
storage[348] = 0;
storage[349] = 0;
storage[350] = 0;
storage[351] = 0;
storage[352] = 0;
storage[353] = 0;
storage[354] = 0;
storage[355] = 0;
storage[356] = 0;
storage[357] = 0;
storage[358] = 0;
storage[359] = 0;
storage[360] = 0;
storage[361] = 0;
storage[362] = 0;
storage[363] = 0;
storage[364] = 0;
storage[365] = 0;
storage[366] = 0;
storage[367] = 0;
storage[368] = 0;
storage[369] = 0;
storage[370] = 0;
storage[371] = 0;
storage[372] = 0;
storage[373] = 0;
storage[374] = 0;
storage[375] = 0;
storage[376] = 0;
storage[377] = 0;
storage[378] = 0;
storage[379] = 0;
storage[380] = 0;
storage[381] = 0;
storage[382] = 0;
storage[383] = 0;
storage[384] = 0;
storage[385] = 0;
storage[386] = 0;
storage[387] = 0;
storage[388] = 0;
storage[389] = 0;
storage[390] = 0;
storage[391] = 0;
storage[392] = 0;
storage[393] = 0;
storage[394] = 0;
storage[395] = 0;
storage[396] = 0;
storage[397] = 0;
storage[398] = 0;
storage[399] = 0;
storage[400] = 0;
storage[401] = 0;
storage[402] = 0;
storage[403] = 0;
storage[404] = 0;
storage[405] = 0;
storage[406] = 0;
storage[407] = 0;
storage[408] = 0;
storage[409] = 0;
storage[410] = 0;
storage[411] = 0;
storage[412] = 0;
storage[413] = 0;
storage[414] = 0;
storage[415] = 0;
storage[416] = 0;
storage[417] = 0;
storage[418] = 0;
storage[419] = 0;
storage[420] = 0;
storage[421] = 0;
storage[422] = 0;
storage[423] = 0;
storage[424] = 0;
storage[425] = 0;
storage[426] = 0;
storage[427] = 0;
storage[428] = 0;
storage[429] = 0;
storage[430] = 0;
storage[431] = 0;
storage[432] = 0;
storage[433] = 0;
storage[434] = 0;
storage[435] = 0;
storage[436] = 0;
storage[437] = 0;
storage[438] = 0;
storage[439] = 0;
storage[440] = 0;
storage[441] = 0;
storage[442] = 0;
storage[443] = 0;
storage[444] = 0;
storage[445] = 0;
storage[446] = 0;
storage[447] = 0;
storage[448] = 0;
storage[449] = 0;
storage[450] = 0;
storage[451] = 0;
storage[452] = 0;
storage[453] = 0;
storage[454] = 0;
storage[455] = 0;
storage[456] = 0;
storage[457] = 0;
storage[458] = 0;
storage[459] = 0;
storage[460] = 0;
storage[461] = 0;
storage[462] = 0;
storage[463] = 0;
storage[464] = 0;
storage[465] = 0;
storage[466] = 0;
storage[467] = 0;
storage[468] = 0;
storage[469] = 0;
storage[470] = 0;
storage[471] = 0;
storage[472] = 0;
storage[473] = 0;
storage[474] = 0;
storage[475] = 0;
storage[476] = 0;
storage[477] = 0;
storage[478] = 0;
storage[479] = 0;
storage[480] = 0;
storage[481] = 0;
storage[482] = 0;
storage[483] = 0;
storage[484] = 0;
storage[485] = 0;
storage[486] = 0;
storage[487] = 0;
storage[488] = 0;
storage[489] = 0;
storage[490] = 0;
storage[491] = 0;
storage[492] = 0;
storage[493] = 0;
storage[494] = 0;
storage[495] = 0;
storage[496] = 0;
storage[497] = 0;
storage[498] = 0;
storage[499] = 0;
storage[500] = 0;
storage[501] = 0;
storage[502] = 0;
storage[503] = 0;
storage[504] = 0;
storage[505] = 0;
storage[506] = 0;
storage[507] = 0;
storage[508] = 0;
storage[509] = 0;
storage[510] = 0;
storage[511] = 0;
storage[512] = 0;
storage[513] = 0;
storage[514] = 0;
storage[515] = 0;
storage[516] = 0;
storage[517] = 0;
storage[518] = 0;
storage[519] = 0;
storage[520] = 0;
storage[521] = 0;
storage[522] = 0;
storage[523] = 0;
storage[524] = 0;
storage[525] = 0;
storage[526] = 0;
storage[527] = 0;
storage[528] = 0;
storage[529] = 0;
storage[530] = 0;
storage[531] = 0;
storage[532] = 0;
storage[533] = 0;
storage[534] = 0;
storage[535] = 0;
storage[536] = 0;
storage[537] = 0;
storage[538] = 0;
storage[539] = 0;
storage[540] = 0;
storage[541] = 0;
storage[542] = 0;
storage[543] = 0;
storage[544] = 0;
storage[545] = 0;
storage[546] = 0;
storage[547] = 0;
storage[548] = 0;
storage[549] = 0;
storage[550] = 0;
storage[551] = 0;
storage[552] = 0;
storage[553] = 0;
storage[554] = 0;
storage[555] = 0;
storage[556] = 0;
storage[557] = 0;
storage[558] = 0;
storage[559] = 0;
storage[560] = 0;
storage[561] = 0;
storage[562] = 0;
storage[563] = 0;
storage[564] = 0;
storage[565] = 0;
storage[566] = 0;
storage[567] = 0;
storage[568] = 0;
storage[569] = 0;
storage[570] = 0;
storage[571] = 0;
storage[572] = 0;
storage[573] = 0;
storage[574] = 0;
storage[575] = 0;
storage[576] = 0;
storage[577] = 0;
storage[578] = 0;
storage[579] = 0;
storage[580] = 0;
storage[581] = 0;
storage[582] = 0;
storage[583] = 0;
storage[584] = 0;
storage[585] = 0;
storage[586] = 0;
storage[587] = 0;
storage[588] = 0;
storage[589] = 0;
storage[590] = 0;
storage[591] = 0;
storage[592] = 0;
storage[593] = 0;
storage[594] = 0;
storage[595] = 0;
storage[596] = 0;
storage[597] = 0;
storage[598] = 0;
storage[599] = 0;
storage[600] = 0;
storage[601] = 0;
storage[602] = 0;
storage[603] = 0;
storage[604] = 0;
storage[605] = 0;
storage[606] = 0;
storage[607] = 0;
storage[608] = 0;
storage[609] = 0;
storage[610] = 0;
storage[611] = 0;
storage[612] = 0;
storage[613] = 0;
storage[614] = 0;
storage[615] = 0;
storage[616] = 0;
storage[617] = 0;
storage[618] = 0;
storage[619] = 0;
storage[620] = 0;
storage[621] = 0;
storage[622] = 0;
storage[623] = 0;
storage[624] = 0;
storage[625] = 0;
storage[626] = 0;
storage[627] = 0;
storage[628] = 0;
storage[629] = 0;
storage[630] = 0;
storage[631] = 0;
storage[632] = 0;
storage[633] = 0;
storage[634] = 0;
storage[635] = 0;
storage[636] = 0;
storage[637] = 0;
storage[638] = 0;
storage[639] = 0;
storage[640] = 0;
storage[641] = 0;
storage[642] = 0;
storage[643] = 0;
storage[644] = 0;
storage[645] = 0;
storage[646] = 0;
storage[647] = 0;
storage[648] = 0;
storage[649] = 0;
storage[650] = 0;
storage[651] = 0;
storage[652] = 0;
storage[653] = 0;
storage[654] = 0;
storage[655] = 0;
storage[656] = 0;
storage[657] = 0;
storage[658] = 0;
storage[659] = 0;
storage[660] = 0;
storage[661] = 0;
storage[662] = 0;
storage[663] = 0;
storage[664] = 0;
storage[665] = 0;
storage[666] = 0;
storage[667] = 0;
storage[668] = 0;
storage[669] = 0;
storage[670] = 0;
storage[671] = 0;
storage[672] = 0;
storage[673] = 0;
storage[674] = 0;
storage[675] = 0;
storage[676] = 0;
storage[677] = 0;
storage[678] = 0;
storage[679] = 0;
storage[680] = 0;
storage[681] = 0;
storage[682] = 0;
storage[683] = 0;
storage[684] = 0;
storage[685] = 0;
storage[686] = 0;
storage[687] = 0;
storage[688] = 0;
storage[689] = 0;
storage[690] = 0;
storage[691] = 0;
storage[692] = 0;
storage[693] = 0;
storage[694] = 0;
storage[695] = 0;
storage[696] = 0;
storage[697] = 0;
storage[698] = 0;
storage[699] = 0;
storage[700] = 0;
storage[701] = 0;
storage[702] = 0;
storage[703] = 0;
storage[704] = 0;
storage[705] = 0;
storage[706] = 0;
storage[707] = 0;
storage[708] = 0;
storage[709] = 0;
storage[710] = 0;
storage[711] = 0;
storage[712] = 0;
storage[713] = 0;
storage[714] = 0;
storage[715] = 0;
storage[716] = 0;
storage[717] = 0;
storage[718] = 0;
storage[719] = 0;
storage[720] = 0;
storage[721] = 0;
storage[722] = 0;
storage[723] = 0;
storage[724] = 0;
storage[725] = 0;
storage[726] = 0;
storage[727] = 0;
storage[728] = 0;
storage[729] = 0;
storage[730] = 0;
storage[731] = 0;
storage[732] = 0;
storage[733] = 0;
storage[734] = 0;
storage[735] = 0;
storage[736] = 0;
storage[737] = 0;
storage[738] = 0;
storage[739] = 0;
storage[740] = 0;
storage[741] = 0;
storage[742] = 0;
storage[743] = 0;
storage[744] = 0;
storage[745] = 0;
storage[746] = 0;
storage[747] = 0;
storage[748] = 0;
storage[749] = 0;
storage[750] = 0;
storage[751] = 0;
storage[752] = 0;
storage[753] = 0;
storage[754] = 0;
storage[755] = 0;
storage[756] = 0;
storage[757] = 0;
storage[758] = 0;
storage[759] = 0;
storage[760] = 0;
storage[761] = 0;
storage[762] = 0;
storage[763] = 0;
storage[764] = 0;
storage[765] = 0;
storage[766] = 0;
storage[767] = 0;
storage[768] = 0;
storage[769] = 0;
storage[770] = 0;
storage[771] = 0;
storage[772] = 0;
storage[773] = 0;
storage[774] = 0;
storage[775] = 0;
storage[776] = 0;
storage[777] = 0;
storage[778] = 0;
storage[779] = 0;
storage[780] = 0;
storage[781] = 0;
storage[782] = 0;
storage[783] = 0;
storage[784] = 0;
storage[785] = 0;
storage[786] = 0;
storage[787] = 0;
storage[788] = 0;
storage[789] = 0;
storage[790] = 0;
storage[791] = 0;
storage[792] = 0;
storage[793] = 0;
storage[794] = 0;
storage[795] = 0;
storage[796] = 0;
storage[797] = 0;
storage[798] = 0;
storage[799] = 0;
storage[800] = 0;
storage[801] = 0;
storage[802] = 0;
storage[803] = 0;
storage[804] = 0;
storage[805] = 0;
storage[806] = 0;
storage[807] = 0;
storage[808] = 0;
storage[809] = 0;
storage[810] = 0;
storage[811] = 0;
storage[812] = 0;
storage[813] = 0;
storage[814] = 0;
storage[815] = 0;
storage[816] = 0;
storage[817] = 0;
storage[818] = 0;
storage[819] = 0;
storage[820] = 0;
storage[821] = 0;
storage[822] = 0;
storage[823] = 0;
storage[824] = 0;
storage[825] = 0;
storage[826] = 0;
storage[827] = 0;
storage[828] = 0;
storage[829] = 0;
storage[830] = 0;
storage[831] = 0;
storage[832] = 0;
storage[833] = 0;
storage[834] = 0;
storage[835] = 0;
storage[836] = 0;
storage[837] = 0;
storage[838] = 0;
storage[839] = 0;
storage[840] = 0;
storage[841] = 0;
storage[842] = 0;
storage[843] = 0;
storage[844] = 0;
storage[845] = 0;
storage[846] = 0;
storage[847] = 0;
storage[848] = 0;
storage[849] = 0;
storage[850] = 0;
storage[851] = 0;
storage[852] = 0;
storage[853] = 0;
storage[854] = 0;
storage[855] = 0;
storage[856] = 0;
storage[857] = 0;
storage[858] = 0;
storage[859] = 0;
storage[860] = 0;
storage[861] = 0;
storage[862] = 0;
storage[863] = 0;
storage[864] = 0;
storage[865] = 0;
storage[866] = 0;
storage[867] = 0;
storage[868] = 0;
storage[869] = 0;
storage[870] = 0;
storage[871] = 0;
storage[872] = 0;
storage[873] = 0;
storage[874] = 0;
storage[875] = 0;
storage[876] = 0;
storage[877] = 0;
storage[878] = 0;
storage[879] = 0;
storage[880] = 0;
storage[881] = 0;
storage[882] = 0;
storage[883] = 0;
storage[884] = 0;
storage[885] = 0;
storage[886] = 0;
storage[887] = 0;
storage[888] = 0;
storage[889] = 0;
storage[890] = 0;
storage[891] = 0;
storage[892] = 0;
storage[893] = 0;
storage[894] = 0;
storage[895] = 0;
storage[896] = 0;
storage[897] = 0;
storage[898] = 0;
storage[899] = 0;
storage[900] = 0;
storage[901] = 0;
storage[902] = 0;
storage[903] = 0;
storage[904] = 0;
storage[905] = 0;
storage[906] = 0;
storage[907] = 0;
storage[908] = 0;
storage[909] = 0;
storage[910] = 0;
storage[911] = 0;
storage[912] = 0;
storage[913] = 0;
storage[914] = 0;
storage[915] = 0;
storage[916] = 0;
storage[917] = 0;
storage[918] = 0;
storage[919] = 0;
storage[920] = 0;
storage[921] = 0;
storage[922] = 0;
storage[923] = 0;
storage[924] = 0;
storage[925] = 0;
storage[926] = 0;
storage[927] = 0;
storage[928] = 0;
storage[929] = 0;
storage[930] = 0;
storage[931] = 0;
storage[932] = 0;
storage[933] = 0;
storage[934] = 0;
storage[935] = 0;
storage[936] = 0;
storage[937] = 0;
storage[938] = 0;
storage[939] = 0;
storage[940] = 0;
storage[941] = 0;
storage[942] = 0;
storage[943] = 0;
storage[944] = 0;
storage[945] = 0;
storage[946] = 0;
storage[947] = 0;
storage[948] = 0;
storage[949] = 0;
storage[950] = 0;
storage[951] = 0;
storage[952] = 0;
storage[953] = 0;
storage[954] = 0;
storage[955] = 0;
storage[956] = 0;
storage[957] = 0;
storage[958] = 0;
storage[959] = 0;
storage[960] = 0;
storage[961] = 0;
storage[962] = 0;
storage[963] = 0;
storage[964] = 0;
storage[965] = 0;
storage[966] = 0;
storage[967] = 0;
storage[968] = 0;
storage[969] = 0;
storage[970] = 0;
storage[971] = 0;
storage[972] = 0;
storage[973] = 0;
storage[974] = 0;
storage[975] = 0;
storage[976] = 0;
storage[977] = 0;
storage[978] = 0;
storage[979] = 0;
storage[980] = 0;
storage[981] = 0;
storage[982] = 0;
storage[983] = 0;
storage[984] = 0;
storage[985] = 0;
storage[986] = 0;
storage[987] = 0;
storage[988] = 0;
storage[989] = 0;
storage[990] = 0;
storage[991] = 0;
storage[992] = 0;
storage[993] = 0;
storage[994] = 0;
storage[995] = 0;
storage[996] = 0;
storage[997] = 0;
storage[998] = 0;
storage[999] = 0;
storage[1000] = 0;
storage[1001] = 0;
storage[1002] = 0;
storage[1003] = 0;
storage[1004] = 0;
storage[1005] = 0;
storage[1006] = 0;
storage[1007] = 0;
storage[1008] = 0;
storage[1009] = 0;
storage[1010] = 0;
storage[1011] = 0;
storage[1012] = 0;
storage[1013] = 0;
storage[1014] = 0;
storage[1015] = 0;
storage[1016] = 0;
storage[1017] = 0;
storage[1018] = 0;
storage[1019] = 0;
storage[1020] = 0;
storage[1021] = 0;
storage[1022] = 0;
storage[1023] = 0;
storage[1024] = 0;
storage[1025] = 0;
storage[1026] = 0;
storage[1027] = 0;
storage[1028] = 0;
storage[1029] = 0;
storage[1030] = 0;
storage[1031] = 0;
storage[1032] = 0;
storage[1033] = 0;
storage[1034] = 0;
storage[1035] = 0;
storage[1036] = 0;
storage[1037] = 0;
storage[1038] = 0;
storage[1039] = 0;
storage[1040] = 0;
storage[1041] = 0;
storage[1042] = 0;
storage[1043] = 0;
storage[1044] = 0;
storage[1045] = 0;
storage[1046] = 0;
storage[1047] = 0;
storage[1048] = 0;
storage[1049] = 0;
storage[1050] = 0;
storage[1051] = 0;
storage[1052] = 0;
storage[1053] = 0;
storage[1054] = 0;
storage[1055] = 0;
storage[1056] = 0;
storage[1057] = 0;
storage[1058] = 0;
storage[1059] = 0;
storage[1060] = 0;
storage[1061] = 0;
storage[1062] = 0;
storage[1063] = 0;
storage[1064] = 0;
storage[1065] = 0;
storage[1066] = 0;
storage[1067] = 0;
storage[1068] = 0;
storage[1069] = 0;
storage[1070] = 0;
storage[1071] = 0;
storage[1072] = 0;
storage[1073] = 0;
storage[1074] = 0;
storage[1075] = 0;
storage[1076] = 0;
storage[1077] = 0;
storage[1078] = 0;
storage[1079] = 0;
storage[1080] = 0;
storage[1081] = 0;
storage[1082] = 0;
storage[1083] = 0;
storage[1084] = 0;
storage[1085] = 0;
storage[1086] = 0;
storage[1087] = 0;
storage[1088] = 0;
storage[1089] = 0;
storage[1090] = 0;
storage[1091] = 0;
storage[1092] = 0;
storage[1093] = 0;
storage[1094] = 0;
storage[1095] = 0;
storage[1096] = 0;
storage[1097] = 0;
storage[1098] = 0;
storage[1099] = 0;
storage[1100] = 0;
storage[1101] = 0;
storage[1102] = 0;
storage[1103] = 0;
storage[1104] = 0;
storage[1105] = 0;
storage[1106] = 0;
storage[1107] = 0;
storage[1108] = 0;
storage[1109] = 0;
storage[1110] = 0;
storage[1111] = 0;
storage[1112] = 0;
storage[1113] = 0;
storage[1114] = 0;
storage[1115] = 0;
storage[1116] = 0;
storage[1117] = 0;
storage[1118] = 0;
storage[1119] = 0;
storage[1120] = 0;
storage[1121] = 0;
storage[1122] = 0;
storage[1123] = 0;
storage[1124] = 0;
storage[1125] = 0;
storage[1126] = 0;
storage[1127] = 0;
storage[1128] = 0;
storage[1129] = 0;
storage[1130] = 0;
storage[1131] = 0;
storage[1132] = 0;
storage[1133] = 0;
storage[1134] = 0;
storage[1135] = 0;
storage[1136] = 0;
storage[1137] = 0;
storage[1138] = 0;
storage[1139] = 0;
storage[1140] = 0;
storage[1141] = 0;
storage[1142] = 0;
storage[1143] = 0;
storage[1144] = 0;
storage[1145] = 0;
storage[1146] = 0;
storage[1147] = 0;
storage[1148] = 0;
storage[1149] = 0;
storage[1150] = 0;
storage[1151] = 0;
storage[1152] = 0;
storage[1153] = 0;
storage[1154] = 0;
storage[1155] = 0;
storage[1156] = 0;
storage[1157] = 0;
storage[1158] = 0;
storage[1159] = 0;
storage[1160] = 0;
storage[1161] = 0;
storage[1162] = 0;
storage[1163] = 0;
storage[1164] = 0;
storage[1165] = 0;
storage[1166] = 0;
storage[1167] = 0;
storage[1168] = 0;
storage[1169] = 0;
storage[1170] = 0;
storage[1171] = 0;
storage[1172] = 0;
storage[1173] = 0;
storage[1174] = 0;
storage[1175] = 0;
storage[1176] = 0;
storage[1177] = 0;
storage[1178] = 0;
storage[1179] = 0;
storage[1180] = 0;
storage[1181] = 0;
storage[1182] = 0;
storage[1183] = 0;
storage[1184] = 0;
storage[1185] = 0;
storage[1186] = 0;
storage[1187] = 0;
storage[1188] = 0;
storage[1189] = 0;
storage[1190] = 0;
storage[1191] = 0;
storage[1192] = 0;
storage[1193] = 0;
storage[1194] = 0;
storage[1195] = 0;
storage[1196] = 0;
storage[1197] = 0;
storage[1198] = 0;
storage[1199] = 0;
storage[1200] = 0;
storage[1201] = 0;
storage[1202] = 0;
storage[1203] = 0;
storage[1204] = 0;
storage[1205] = 0;
storage[1206] = 0;
storage[1207] = 0;
storage[1208] = 0;
storage[1209] = 0;
storage[1210] = 0;
storage[1211] = 0;
storage[1212] = 0;
storage[1213] = 0;
storage[1214] = 0;
storage[1215] = 0;
storage[1216] = 0;
storage[1217] = 0;
storage[1218] = 0;
storage[1219] = 0;
storage[1220] = 0;
storage[1221] = 0;
storage[1222] = 0;
storage[1223] = 0;
storage[1224] = 0;
storage[1225] = 0;
storage[1226] = 0;
storage[1227] = 0;
storage[1228] = 0;
storage[1229] = 0;
storage[1230] = 0;
storage[1231] = 0;
storage[1232] = 0;
storage[1233] = 0;
storage[1234] = 0;
storage[1235] = 0;
storage[1236] = 0;
storage[1237] = 0;
storage[1238] = 0;
storage[1239] = 0;
storage[1240] = 0;
storage[1241] = 0;
storage[1242] = 0;
storage[1243] = 0;
storage[1244] = 0;
storage[1245] = 0;
storage[1246] = 0;
storage[1247] = 0;
storage[1248] = 0;
storage[1249] = 0;
storage[1250] = 0;
storage[1251] = 0;
storage[1252] = 0;
storage[1253] = 0;
storage[1254] = 0;
storage[1255] = 0;
storage[1256] = 0;
storage[1257] = 0;
storage[1258] = 0;
storage[1259] = 0;
storage[1260] = 0;
storage[1261] = 0;
storage[1262] = 0;
storage[1263] = 0;
storage[1264] = 0;
storage[1265] = 0;
storage[1266] = 0;
storage[1267] = 0;
storage[1268] = 0;
storage[1269] = 0;
storage[1270] = 0;
storage[1271] = 0;
storage[1272] = 0;
storage[1273] = 0;
storage[1274] = 0;
storage[1275] = 0;
storage[1276] = 0;
storage[1277] = 0;
storage[1278] = 0;
storage[1279] = 0;
storage[1280] = 0;
storage[1281] = 0;
storage[1282] = 0;
storage[1283] = 0;
storage[1284] = 0;
storage[1285] = 0;
storage[1286] = 0;
storage[1287] = 0;
storage[1288] = 0;
storage[1289] = 0;
storage[1290] = 0;
storage[1291] = 0;
storage[1292] = 0;
storage[1293] = 0;
storage[1294] = 0;
storage[1295] = 0;
storage[1296] = 0;
storage[1297] = 0;
storage[1298] = 0;
storage[1299] = 0;
storage[1300] = 0;
storage[1301] = 0;
storage[1302] = 0;
storage[1303] = 0;
storage[1304] = 0;
storage[1305] = 0;
storage[1306] = 0;
storage[1307] = 0;
storage[1308] = 0;
storage[1309] = 0;
storage[1310] = 0;
storage[1311] = 0;
storage[1312] = 0;
storage[1313] = 0;
storage[1314] = 0;
storage[1315] = 0;
storage[1316] = 0;
storage[1317] = 0;
storage[1318] = 0;
storage[1319] = 0;
storage[1320] = 0;
storage[1321] = 0;
storage[1322] = 0;
storage[1323] = 0;
storage[1324] = 0;
storage[1325] = 0;
storage[1326] = 0;
storage[1327] = 0;
storage[1328] = 0;
storage[1329] = 0;
storage[1330] = 0;
storage[1331] = 0;
storage[1332] = 0;
storage[1333] = 0;
storage[1334] = 0;
storage[1335] = 0;
storage[1336] = 0;
storage[1337] = 0;
storage[1338] = 0;
storage[1339] = 0;
storage[1340] = 0;
storage[1341] = 0;
storage[1342] = 0;
storage[1343] = 0;
storage[1344] = 0;
storage[1345] = 0;
storage[1346] = 0;
storage[1347] = 0;
storage[1348] = 0;
storage[1349] = 0;
storage[1350] = 0;
storage[1351] = 0;
storage[1352] = 0;
storage[1353] = 0;
storage[1354] = 0;
storage[1355] = 0;
storage[1356] = 0;
storage[1357] = 0;
storage[1358] = 0;
storage[1359] = 0;
storage[1360] = 0;
storage[1361] = 0;
storage[1362] = 0;
storage[1363] = 0;
storage[1364] = 0;
storage[1365] = 0;
storage[1366] = 0;
storage[1367] = 0;
storage[1368] = 0;
storage[1369] = 0;
storage[1370] = 0;
storage[1371] = 0;
storage[1372] = 0;
storage[1373] = 0;
storage[1374] = 0;
storage[1375] = 0;
storage[1376] = 0;
storage[1377] = 0;
storage[1378] = 0;
storage[1379] = 0;
storage[1380] = 0;
storage[1381] = 0;
storage[1382] = 0;
storage[1383] = 0;
storage[1384] = 0;
storage[1385] = 0;
storage[1386] = 0;
storage[1387] = 0;
storage[1388] = 0;
storage[1389] = 0;
storage[1390] = 0;
storage[1391] = 0;
storage[1392] = 0;
storage[1393] = 0;
storage[1394] = 0;
storage[1395] = 0;
storage[1396] = 0;
storage[1397] = 0;
storage[1398] = 0;
storage[1399] = 0;
storage[1400] = 0;
storage[1401] = 0;
storage[1402] = 0;
storage[1403] = 0;
storage[1404] = 0;
storage[1405] = 0;
storage[1406] = 0;
storage[1407] = 0;
storage[1408] = 0;
storage[1409] = 0;
storage[1410] = 0;
storage[1411] = 0;
storage[1412] = 0;
storage[1413] = 0;
storage[1414] = 0;
storage[1415] = 0;
storage[1416] = 0;
storage[1417] = 0;
storage[1418] = 0;
storage[1419] = 0;
storage[1420] = 0;
storage[1421] = 0;
storage[1422] = 0;
storage[1423] = 0;
storage[1424] = 0;
storage[1425] = 0;
storage[1426] = 0;
storage[1427] = 0;
storage[1428] = 0;
storage[1429] = 0;
storage[1430] = 0;
storage[1431] = 0;
storage[1432] = 0;
storage[1433] = 0;
storage[1434] = 0;
storage[1435] = 0;
storage[1436] = 0;
storage[1437] = 0;
storage[1438] = 0;
storage[1439] = 0;
storage[1440] = 0;
storage[1441] = 0;
storage[1442] = 0;
storage[1443] = 0;
storage[1444] = 0;
storage[1445] = 0;
storage[1446] = 0;
storage[1447] = 0;
storage[1448] = 0;
storage[1449] = 0;
storage[1450] = 0;
storage[1451] = 0;
storage[1452] = 0;
storage[1453] = 0;
storage[1454] = 0;
storage[1455] = 0;
storage[1456] = 0;
storage[1457] = 0;
storage[1458] = 0;
storage[1459] = 0;
storage[1460] = 0;
storage[1461] = 0;
storage[1462] = 0;
storage[1463] = 0;
storage[1464] = 0;
storage[1465] = 0;
storage[1466] = 0;
storage[1467] = 0;
storage[1468] = 0;
storage[1469] = 0;
storage[1470] = 0;
storage[1471] = 0;
storage[1472] = 0;
storage[1473] = 0;
storage[1474] = 0;
storage[1475] = 0;
storage[1476] = 0;
storage[1477] = 0;
storage[1478] = 0;
storage[1479] = 0;
storage[1480] = 0;
storage[1481] = 0;
storage[1482] = 0;
storage[1483] = 0;
storage[1484] = 0;
storage[1485] = 0;
storage[1486] = 0;
storage[1487] = 0;
storage[1488] = 0;
storage[1489] = 0;
storage[1490] = 0;
storage[1491] = 0;
storage[1492] = 0;
storage[1493] = 0;
storage[1494] = 0;
storage[1495] = 0;
storage[1496] = 0;
storage[1497] = 0;
storage[1498] = 0;
storage[1499] = 0;
storage[1500] = 0;
storage[1501] = 0;
storage[1502] = 0;
storage[1503] = 0;
storage[1504] = 0;
storage[1505] = 0;
storage[1506] = 0;
storage[1507] = 0;
storage[1508] = 0;
storage[1509] = 0;
storage[1510] = 0;
storage[1511] = 0;
storage[1512] = 0;
storage[1513] = 0;
storage[1514] = 0;
storage[1515] = 0;
storage[1516] = 0;
storage[1517] = 0;
storage[1518] = 0;
storage[1519] = 0;
storage[1520] = 0;
storage[1521] = 0;
storage[1522] = 0;
storage[1523] = 0;
storage[1524] = 0;
storage[1525] = 0;
storage[1526] = 0;
storage[1527] = 0;
storage[1528] = 0;
storage[1529] = 0;
storage[1530] = 0;
storage[1531] = 0;
storage[1532] = 0;
storage[1533] = 0;
storage[1534] = 0;
storage[1535] = 0;
storage[1536] = 0;
storage[1537] = 0;
storage[1538] = 0;
storage[1539] = 0;
storage[1540] = 0;
storage[1541] = 0;
storage[1542] = 0;
storage[1543] = 0;
storage[1544] = 0;
storage[1545] = 0;
storage[1546] = 0;
storage[1547] = 0;
storage[1548] = 0;
storage[1549] = 0;
storage[1550] = 0;
storage[1551] = 0;
storage[1552] = 0;
storage[1553] = 0;
storage[1554] = 0;
storage[1555] = 0;
storage[1556] = 0;
storage[1557] = 0;
storage[1558] = 0;
storage[1559] = 0;
storage[1560] = 0;
storage[1561] = 0;
storage[1562] = 0;
storage[1563] = 0;
storage[1564] = 0;
storage[1565] = 0;
storage[1566] = 0;
storage[1567] = 0;
storage[1568] = 0;
storage[1569] = 0;
storage[1570] = 0;
storage[1571] = 0;
storage[1572] = 0;
storage[1573] = 0;
storage[1574] = 0;
storage[1575] = 0;
storage[1576] = 0;
storage[1577] = 0;
storage[1578] = 0;
storage[1579] = 0;
storage[1580] = 0;
storage[1581] = 0;
storage[1582] = 0;
storage[1583] = 0;
storage[1584] = 0;
storage[1585] = 0;
storage[1586] = 0;
storage[1587] = 0;
storage[1588] = 0;
storage[1589] = 0;
storage[1590] = 0;
storage[1591] = 0;
storage[1592] = 0;
storage[1593] = 0;
storage[1594] = 0;
storage[1595] = 0;
storage[1596] = 0;
storage[1597] = 0;
storage[1598] = 0;
storage[1599] = 0;
storage[1600] = 0;
storage[1601] = 0;
storage[1602] = 0;
storage[1603] = 0;
storage[1604] = 0;
storage[1605] = 0;
storage[1606] = 0;
storage[1607] = 0;
storage[1608] = 0;
storage[1609] = 0;
storage[1610] = 0;
storage[1611] = 0;
storage[1612] = 0;
storage[1613] = 0;
storage[1614] = 0;
storage[1615] = 0;
storage[1616] = 0;
storage[1617] = 0;
storage[1618] = 0;
storage[1619] = 0;
storage[1620] = 0;
storage[1621] = 0;
storage[1622] = 0;
storage[1623] = 0;
storage[1624] = 0;
storage[1625] = 0;
storage[1626] = 0;
storage[1627] = 0;
storage[1628] = 0;
storage[1629] = 0;
storage[1630] = 0;
storage[1631] = 0;
storage[1632] = 0;
storage[1633] = 0;
storage[1634] = 0;
storage[1635] = 0;
storage[1636] = 0;
storage[1637] = 0;
storage[1638] = 0;
storage[1639] = 0;
storage[1640] = 0;
storage[1641] = 0;
storage[1642] = 0;
storage[1643] = 0;
storage[1644] = 0;
storage[1645] = 0;
storage[1646] = 0;
storage[1647] = 0;
storage[1648] = 0;
storage[1649] = 0;
storage[1650] = 0;
storage[1651] = 0;
storage[1652] = 0;
storage[1653] = 0;
storage[1654] = 0;
storage[1655] = 0;
storage[1656] = 0;
storage[1657] = 0;
storage[1658] = 0;
storage[1659] = 0;
storage[1660] = 0;
storage[1661] = 0;
storage[1662] = 0;
storage[1663] = 0;
storage[1664] = 0;
storage[1665] = 0;
storage[1666] = 0;
storage[1667] = 0;
storage[1668] = 0;
storage[1669] = 0;
storage[1670] = 0;
storage[1671] = 0;
storage[1672] = 0;
storage[1673] = 0;
storage[1674] = 0;
storage[1675] = 0;
storage[1676] = 0;
storage[1677] = 0;
storage[1678] = 0;
storage[1679] = 0;
storage[1680] = 0;
storage[1681] = 0;
storage[1682] = 0;
storage[1683] = 0;
storage[1684] = 0;
storage[1685] = 0;
storage[1686] = 0;
storage[1687] = 0;
storage[1688] = 0;
storage[1689] = 0;
storage[1690] = 0;
storage[1691] = 0;
storage[1692] = 0;
storage[1693] = 0;
storage[1694] = 0;
storage[1695] = 0;
storage[1696] = 0;
storage[1697] = 0;
storage[1698] = 0;
storage[1699] = 0;
storage[1700] = 0;
storage[1701] = 0;
storage[1702] = 0;
storage[1703] = 0;
storage[1704] = 0;
storage[1705] = 0;
storage[1706] = 0;
storage[1707] = 0;
storage[1708] = 0;
storage[1709] = 0;
storage[1710] = 0;
storage[1711] = 0;
storage[1712] = 0;
storage[1713] = 0;
storage[1714] = 0;
storage[1715] = 0;
storage[1716] = 0;
storage[1717] = 0;
storage[1718] = 0;
storage[1719] = 0;
storage[1720] = 0;
storage[1721] = 0;
storage[1722] = 0;
storage[1723] = 0;
storage[1724] = 0;
storage[1725] = 0;
storage[1726] = 0;
storage[1727] = 0;
storage[1728] = 0;
storage[1729] = 0;
storage[1730] = 0;
storage[1731] = 0;
storage[1732] = 0;
storage[1733] = 0;
storage[1734] = 0;
storage[1735] = 0;
storage[1736] = 0;
storage[1737] = 0;
storage[1738] = 0;
storage[1739] = 0;
storage[1740] = 0;
storage[1741] = 0;
storage[1742] = 0;
storage[1743] = 0;
storage[1744] = 0;
storage[1745] = 0;
storage[1746] = 0;
storage[1747] = 0;
storage[1748] = 0;
storage[1749] = 0;
storage[1750] = 0;
storage[1751] = 0;
storage[1752] = 0;
storage[1753] = 0;
storage[1754] = 0;
storage[1755] = 0;
storage[1756] = 0;
storage[1757] = 0;
storage[1758] = 0;
storage[1759] = 0;
storage[1760] = 0;
storage[1761] = 0;
storage[1762] = 0;
storage[1763] = 0;
storage[1764] = 0;
storage[1765] = 0;
storage[1766] = 0;
storage[1767] = 0;
storage[1768] = 0;
storage[1769] = 0;
storage[1770] = 0;
storage[1771] = 0;
storage[1772] = 0;
storage[1773] = 0;
storage[1774] = 0;
storage[1775] = 0;
storage[1776] = 0;
storage[1777] = 0;
storage[1778] = 0;
storage[1779] = 0;
storage[1780] = 0;
storage[1781] = 0;
storage[1782] = 0;
storage[1783] = 0;
storage[1784] = 0;
storage[1785] = 0;
storage[1786] = 0;
storage[1787] = 0;
storage[1788] = 0;
storage[1789] = 0;
storage[1790] = 0;
storage[1791] = 0;
storage[1792] = 0;
storage[1793] = 0;
storage[1794] = 0;
storage[1795] = 0;
storage[1796] = 0;
storage[1797] = 0;
storage[1798] = 0;
storage[1799] = 0;
storage[1800] = 0;
storage[1801] = 0;
storage[1802] = 0;
storage[1803] = 0;
storage[1804] = 0;
storage[1805] = 0;
storage[1806] = 0;
storage[1807] = 0;
storage[1808] = 0;
storage[1809] = 0;
storage[1810] = 0;
storage[1811] = 0;
storage[1812] = 0;
storage[1813] = 0;
storage[1814] = 0;
storage[1815] = 0;
storage[1816] = 0;
storage[1817] = 0;
storage[1818] = 0;
storage[1819] = 0;
storage[1820] = 0;
storage[1821] = 0;
storage[1822] = 0;
storage[1823] = 0;
storage[1824] = 0;
storage[1825] = 0;
storage[1826] = 0;
storage[1827] = 0;
storage[1828] = 0;
storage[1829] = 0;
storage[1830] = 0;
storage[1831] = 0;
storage[1832] = 0;
storage[1833] = 0;
storage[1834] = 0;
storage[1835] = 0;
storage[1836] = 0;
storage[1837] = 0;
storage[1838] = 0;
storage[1839] = 0;
storage[1840] = 0;
storage[1841] = 0;
storage[1842] = 0;
storage[1843] = 0;
storage[1844] = 0;
storage[1845] = 0;
storage[1846] = 0;
storage[1847] = 0;
storage[1848] = 0;
storage[1849] = 0;
storage[1850] = 0;
storage[1851] = 0;
storage[1852] = 0;
storage[1853] = 0;
storage[1854] = 0;
storage[1855] = 0;
storage[1856] = 0;
storage[1857] = 0;
storage[1858] = 0;
storage[1859] = 0;
storage[1860] = 0;
storage[1861] = 0;
storage[1862] = 0;
storage[1863] = 0;
storage[1864] = 0;
storage[1865] = 0;
storage[1866] = 0;
storage[1867] = 0;
storage[1868] = 0;
storage[1869] = 0;
storage[1870] = 0;
storage[1871] = 0;
storage[1872] = 0;
storage[1873] = 0;
storage[1874] = 0;
storage[1875] = 0;
storage[1876] = 0;
storage[1877] = 0;
storage[1878] = 0;
storage[1879] = 0;
storage[1880] = 0;
storage[1881] = 0;
storage[1882] = 0;
storage[1883] = 0;
storage[1884] = 0;
storage[1885] = 0;
storage[1886] = 0;
storage[1887] = 0;
storage[1888] = 0;
storage[1889] = 0;
storage[1890] = 0;
storage[1891] = 0;
storage[1892] = 0;
storage[1893] = 0;
storage[1894] = 0;
storage[1895] = 0;
storage[1896] = 0;
storage[1897] = 0;
storage[1898] = 0;
storage[1899] = 0;
storage[1900] = 0;
storage[1901] = 0;
storage[1902] = 0;
storage[1903] = 0;
storage[1904] = 0;
storage[1905] = 0;
storage[1906] = 0;
storage[1907] = 0;
storage[1908] = 0;
storage[1909] = 0;
storage[1910] = 0;
storage[1911] = 0;
storage[1912] = 0;
storage[1913] = 0;
storage[1914] = 0;
storage[1915] = 0;
storage[1916] = 0;
storage[1917] = 0;
storage[1918] = 0;
storage[1919] = 0;
storage[1920] = 0;
storage[1921] = 0;
storage[1922] = 0;
storage[1923] = 0;
storage[1924] = 0;
storage[1925] = 0;
storage[1926] = 0;
storage[1927] = 0;
storage[1928] = 0;
storage[1929] = 0;
storage[1930] = 0;
storage[1931] = 0;
storage[1932] = 0;
storage[1933] = 0;
storage[1934] = 0;
storage[1935] = 0;
storage[1936] = 0;
storage[1937] = 0;
storage[1938] = 0;
storage[1939] = 0;
storage[1940] = 0;
storage[1941] = 0;
storage[1942] = 0;
storage[1943] = 0;
storage[1944] = 0;
storage[1945] = 0;
storage[1946] = 0;
storage[1947] = 0;
storage[1948] = 0;
storage[1949] = 0;
storage[1950] = 0;
storage[1951] = 0;
storage[1952] = 0;
storage[1953] = 0;
storage[1954] = 0;
storage[1955] = 0;
storage[1956] = 0;
storage[1957] = 0;
storage[1958] = 0;
storage[1959] = 0;
storage[1960] = 0;
storage[1961] = 0;
storage[1962] = 0;
storage[1963] = 0;
storage[1964] = 0;
storage[1965] = 0;
storage[1966] = 0;
storage[1967] = 0;
storage[1968] = 0;
storage[1969] = 0;
storage[1970] = 0;
storage[1971] = 0;
storage[1972] = 0;
storage[1973] = 0;
storage[1974] = 0;
storage[1975] = 0;
storage[1976] = 0;
storage[1977] = 0;
storage[1978] = 0;
storage[1979] = 0;
storage[1980] = 0;
storage[1981] = 0;
storage[1982] = 0;
storage[1983] = 0;
storage[1984] = 0;
storage[1985] = 0;
storage[1986] = 0;
storage[1987] = 0;
storage[1988] = 0;
storage[1989] = 0;
storage[1990] = 0;
storage[1991] = 0;
storage[1992] = 0;
storage[1993] = 0;
storage[1994] = 0;
storage[1995] = 0;
storage[1996] = 0;
storage[1997] = 0;
storage[1998] = 0;
storage[1999] = 0;
storage[2000] = 0;
storage[2001] = 0;
storage[2002] = 0;
storage[2003] = 0;
storage[2004] = 0;
storage[2005] = 0;
storage[2006] = 0;
storage[2007] = 0;
storage[2008] = 0;
storage[2009] = 0;
storage[2010] = 0;
storage[2011] = 0;
storage[2012] = 0;
storage[2013] = 0;
storage[2014] = 0;
storage[2015] = 0;
storage[2016] = 0;
storage[2017] = 0;
storage[2018] = 0;
storage[2019] = 0;
storage[2020] = 0;
storage[2021] = 0;
storage[2022] = 0;
storage[2023] = 0;
storage[2024] = 0;
storage[2025] = 0;
storage[2026] = 0;
storage[2027] = 0;
storage[2028] = 0;
storage[2029] = 0;
storage[2030] = 0;
storage[2031] = 0;
storage[2032] = 0;
storage[2033] = 0;
storage[2034] = 0;
storage[2035] = 0;
storage[2036] = 0;
storage[2037] = 0;
storage[2038] = 0;
storage[2039] = 0;
storage[2040] = 0;
storage[2041] = 0;
storage[2042] = 0;
storage[2043] = 0;
storage[2044] = 0;
storage[2045] = 0;
storage[2046] = 0;
storage[2047] = 0;
storage[2048] = 0;
storage[2049] = 0;
storage[2050] = 0;
storage[2051] = 0;
storage[2052] = 0;
storage[2053] = 0;
storage[2054] = 0;
storage[2055] = 0;
storage[2056] = 0;
storage[2057] = 0;
storage[2058] = 0;
storage[2059] = 0;
storage[2060] = 0;
storage[2061] = 0;
storage[2062] = 0;
storage[2063] = 0;
storage[2064] = 0;
storage[2065] = 0;
storage[2066] = 0;
storage[2067] = 0;
storage[2068] = 0;
storage[2069] = 0;
storage[2070] = 0;
storage[2071] = 0;
storage[2072] = 0;
storage[2073] = 0;
storage[2074] = 0;
storage[2075] = 0;
storage[2076] = 0;
storage[2077] = 0;
storage[2078] = 0;
storage[2079] = 0;
storage[2080] = 0;
storage[2081] = 0;
storage[2082] = 0;
storage[2083] = 0;
storage[2084] = 0;
storage[2085] = 0;
storage[2086] = 0;
storage[2087] = 0;
storage[2088] = 0;
storage[2089] = 0;
storage[2090] = 0;
storage[2091] = 0;
storage[2092] = 0;
storage[2093] = 0;
storage[2094] = 0;
storage[2095] = 0;
storage[2096] = 0;
storage[2097] = 0;
storage[2098] = 0;
storage[2099] = 0;
storage[2100] = 0;
storage[2101] = 0;
storage[2102] = 0;
storage[2103] = 0;
storage[2104] = 0;
storage[2105] = 0;
storage[2106] = 0;
storage[2107] = 0;
storage[2108] = 0;
storage[2109] = 0;
storage[2110] = 0;
storage[2111] = 0;
storage[2112] = 0;
storage[2113] = 0;
storage[2114] = 0;
storage[2115] = 0;
storage[2116] = 0;
storage[2117] = 0;
storage[2118] = 0;
storage[2119] = 0;
storage[2120] = 0;
storage[2121] = 0;
storage[2122] = 0;
storage[2123] = 0;
storage[2124] = 0;
storage[2125] = 0;
storage[2126] = 0;
storage[2127] = 0;
storage[2128] = 0;
storage[2129] = 0;
storage[2130] = 0;
storage[2131] = 0;
storage[2132] = 0;
storage[2133] = 0;
storage[2134] = 0;
storage[2135] = 0;
storage[2136] = 0;
storage[2137] = 0;
storage[2138] = 0;
storage[2139] = 0;
storage[2140] = 0;
storage[2141] = 0;
storage[2142] = 0;
storage[2143] = 0;
storage[2144] = 0;
storage[2145] = 0;
storage[2146] = 0;
storage[2147] = 0;
storage[2148] = 0;
storage[2149] = 0;
storage[2150] = 0;
storage[2151] = 0;
storage[2152] = 0;
storage[2153] = 0;
storage[2154] = 0;
storage[2155] = 0;
storage[2156] = 0;
storage[2157] = 0;
storage[2158] = 0;
storage[2159] = 0;
storage[2160] = 0;
storage[2161] = 0;
storage[2162] = 0;
storage[2163] = 0;
storage[2164] = 0;
storage[2165] = 0;
storage[2166] = 0;
storage[2167] = 0;
storage[2168] = 0;
storage[2169] = 0;
storage[2170] = 0;
storage[2171] = 0;
storage[2172] = 0;
storage[2173] = 0;
storage[2174] = 0;
storage[2175] = 0;
storage[2176] = 0;
storage[2177] = 0;
storage[2178] = 0;
storage[2179] = 0;
storage[2180] = 0;
storage[2181] = 0;
storage[2182] = 0;
storage[2183] = 0;
storage[2184] = 0;
storage[2185] = 0;
storage[2186] = 0;
storage[2187] = 0;
storage[2188] = 0;
storage[2189] = 0;
storage[2190] = 0;
storage[2191] = 0;
storage[2192] = 0;
storage[2193] = 0;
storage[2194] = 0;
storage[2195] = 0;
storage[2196] = 0;
storage[2197] = 0;
storage[2198] = 0;
storage[2199] = 0;
storage[2200] = 0;
storage[2201] = 0;
storage[2202] = 0;
storage[2203] = 0;
storage[2204] = 0;
storage[2205] = 0;
storage[2206] = 0;
storage[2207] = 0;
storage[2208] = 0;
storage[2209] = 0;
storage[2210] = 0;
storage[2211] = 0;
storage[2212] = 0;
storage[2213] = 0;
storage[2214] = 0;
storage[2215] = 0;
storage[2216] = 0;
storage[2217] = 0;
storage[2218] = 0;
storage[2219] = 0;
storage[2220] = 0;
storage[2221] = 0;
storage[2222] = 0;
storage[2223] = 0;
storage[2224] = 0;
storage[2225] = 0;
storage[2226] = 0;
storage[2227] = 0;
storage[2228] = 0;
storage[2229] = 0;
storage[2230] = 0;
storage[2231] = 0;
storage[2232] = 0;
storage[2233] = 0;
storage[2234] = 0;
storage[2235] = 0;
storage[2236] = 0;
storage[2237] = 0;
storage[2238] = 0;
storage[2239] = 0;
storage[2240] = 0;
storage[2241] = 0;
storage[2242] = 0;
storage[2243] = 0;
storage[2244] = 0;
storage[2245] = 0;
storage[2246] = 0;
storage[2247] = 0;
storage[2248] = 0;
storage[2249] = 0;
storage[2250] = 0;
storage[2251] = 0;
storage[2252] = 0;
storage[2253] = 0;
storage[2254] = 0;
storage[2255] = 0;
storage[2256] = 0;
storage[2257] = 0;
storage[2258] = 0;
storage[2259] = 0;
storage[2260] = 0;
storage[2261] = 0;
storage[2262] = 0;
storage[2263] = 0;
storage[2264] = 0;
storage[2265] = 0;
storage[2266] = 0;
storage[2267] = 0;
storage[2268] = 0;
storage[2269] = 0;
storage[2270] = 0;
storage[2271] = 0;
storage[2272] = 0;
storage[2273] = 0;
storage[2274] = 0;
storage[2275] = 0;
storage[2276] = 0;
storage[2277] = 0;
storage[2278] = 0;
storage[2279] = 0;
storage[2280] = 0;
storage[2281] = 0;
storage[2282] = 0;
storage[2283] = 0;
storage[2284] = 0;
storage[2285] = 0;
storage[2286] = 0;
storage[2287] = 0;
storage[2288] = 0;
storage[2289] = 0;
storage[2290] = 0;
storage[2291] = 0;
storage[2292] = 0;
storage[2293] = 0;
storage[2294] = 0;
storage[2295] = 0;
storage[2296] = 0;
storage[2297] = 0;
storage[2298] = 0;
storage[2299] = 0;
storage[2300] = 0;
storage[2301] = 0;
storage[2302] = 0;
storage[2303] = 0;
storage[2304] = 0;
storage[2305] = 0;
storage[2306] = 0;
storage[2307] = 0;
storage[2308] = 0;
storage[2309] = 0;
storage[2310] = 0;
storage[2311] = 0;
storage[2312] = 0;
storage[2313] = 0;
storage[2314] = 0;
storage[2315] = 0;
storage[2316] = 0;
storage[2317] = 0;
storage[2318] = 0;
storage[2319] = 0;
storage[2320] = 0;
storage[2321] = 0;
storage[2322] = 0;
storage[2323] = 0;
storage[2324] = 0;
storage[2325] = 0;
storage[2326] = 0;
storage[2327] = 0;
storage[2328] = 0;
storage[2329] = 0;
storage[2330] = 0;
storage[2331] = 0;
storage[2332] = 0;
storage[2333] = 0;
storage[2334] = 0;
storage[2335] = 0;
storage[2336] = 0;
storage[2337] = 0;
storage[2338] = 0;
storage[2339] = 0;
storage[2340] = 0;
storage[2341] = 0;
storage[2342] = 0;
storage[2343] = 0;
storage[2344] = 0;
storage[2345] = 0;
storage[2346] = 0;
storage[2347] = 0;
storage[2348] = 0;
storage[2349] = 0;
storage[2350] = 0;
storage[2351] = 0;
storage[2352] = 0;
storage[2353] = 0;
storage[2354] = 0;
storage[2355] = 0;
storage[2356] = 0;
storage[2357] = 0;
storage[2358] = 0;
storage[2359] = 0;
storage[2360] = 0;
storage[2361] = 0;
storage[2362] = 0;
storage[2363] = 0;
storage[2364] = 0;
storage[2365] = 0;
storage[2366] = 0;
storage[2367] = 0;
storage[2368] = 0;
storage[2369] = 0;
storage[2370] = 0;
storage[2371] = 0;
storage[2372] = 0;
storage[2373] = 0;
storage[2374] = 0;
storage[2375] = 0;
storage[2376] = 0;
storage[2377] = 0;
storage[2378] = 0;
storage[2379] = 0;
storage[2380] = 0;
storage[2381] = 0;
storage[2382] = 0;
storage[2383] = 0;
storage[2384] = 0;
storage[2385] = 0;
storage[2386] = 0;
storage[2387] = 0;
storage[2388] = 0;
storage[2389] = 0;
storage[2390] = 0;
storage[2391] = 0;
storage[2392] = 0;
storage[2393] = 0;
storage[2394] = 0;
storage[2395] = 0;
storage[2396] = 0;
storage[2397] = 0;
storage[2398] = 0;
storage[2399] = 0;
storage[2400] = 0;
storage[2401] = 0;
storage[2402] = 0;
storage[2403] = 0;
storage[2404] = 0;
storage[2405] = 0;
storage[2406] = 0;
storage[2407] = 0;
storage[2408] = 0;
storage[2409] = 0;
storage[2410] = 0;
storage[2411] = 0;
storage[2412] = 0;
storage[2413] = 0;
storage[2414] = 0;
storage[2415] = 0;
storage[2416] = 0;
storage[2417] = 0;
storage[2418] = 0;
storage[2419] = 0;
storage[2420] = 0;
storage[2421] = 0;
storage[2422] = 0;
storage[2423] = 0;
storage[2424] = 0;
storage[2425] = 0;
storage[2426] = 0;
storage[2427] = 0;
storage[2428] = 0;
storage[2429] = 0;
storage[2430] = 0;
storage[2431] = 0;
storage[2432] = 0;
storage[2433] = 0;
storage[2434] = 0;
storage[2435] = 0;
storage[2436] = 0;
storage[2437] = 0;
storage[2438] = 0;
storage[2439] = 0;
storage[2440] = 0;
storage[2441] = 0;
storage[2442] = 0;
storage[2443] = 0;
storage[2444] = 0;
storage[2445] = 0;
storage[2446] = 0;
storage[2447] = 0;
storage[2448] = 0;
storage[2449] = 0;
storage[2450] = 0;
storage[2451] = 0;
storage[2452] = 0;
storage[2453] = 0;
storage[2454] = 0;
storage[2455] = 0;
storage[2456] = 0;
storage[2457] = 0;
storage[2458] = 0;
storage[2459] = 0;
storage[2460] = 0;
storage[2461] = 0;
storage[2462] = 0;
storage[2463] = 0;
storage[2464] = 0;
storage[2465] = 0;
storage[2466] = 0;
storage[2467] = 0;
storage[2468] = 0;
storage[2469] = 0;
storage[2470] = 0;
storage[2471] = 0;
storage[2472] = 0;
storage[2473] = 0;
storage[2474] = 0;
storage[2475] = 0;
storage[2476] = 0;
storage[2477] = 0;
storage[2478] = 0;
storage[2479] = 0;
storage[2480] = 0;
storage[2481] = 0;
storage[2482] = 0;
storage[2483] = 0;
storage[2484] = 0;
storage[2485] = 0;
storage[2486] = 0;
storage[2487] = 0;
storage[2488] = 0;
storage[2489] = 0;
storage[2490] = 0;
storage[2491] = 0;
storage[2492] = 0;
storage[2493] = 0;
storage[2494] = 0;
storage[2495] = 0;
storage[2496] = 0;
storage[2497] = 0;
storage[2498] = 0;
storage[2499] = 0;
storage[2500] = 0;
storage[2501] = 0;
storage[2502] = 0;
storage[2503] = 0;
storage[2504] = 0;
storage[2505] = 0;
storage[2506] = 0;
storage[2507] = 0;
storage[2508] = 0;
storage[2509] = 0;
storage[2510] = 0;
storage[2511] = 0;
storage[2512] = 0;
storage[2513] = 0;
storage[2514] = 0;
storage[2515] = 0;
storage[2516] = 0;
storage[2517] = 0;
storage[2518] = 0;
storage[2519] = 0;
storage[2520] = 0;
storage[2521] = 0;
storage[2522] = 0;
storage[2523] = 0;
storage[2524] = 0;
storage[2525] = 0;
storage[2526] = 0;
storage[2527] = 0;
storage[2528] = 0;
storage[2529] = 0;
storage[2530] = 0;
storage[2531] = 0;
storage[2532] = 0;
storage[2533] = 0;
storage[2534] = 0;
storage[2535] = 0;
storage[2536] = 0;
storage[2537] = 0;
storage[2538] = 0;
storage[2539] = 0;
storage[2540] = 0;
storage[2541] = 0;
storage[2542] = 0;
storage[2543] = 0;
storage[2544] = 0;
storage[2545] = 0;
storage[2546] = 0;
storage[2547] = 0;
storage[2548] = 0;
storage[2549] = 0;
storage[2550] = 0;
storage[2551] = 0;
storage[2552] = 0;
storage[2553] = 0;
storage[2554] = 0;
storage[2555] = 0;
storage[2556] = 0;
storage[2557] = 0;
storage[2558] = 0;
storage[2559] = 0;
storage[2560] = 0;
storage[2561] = 0;
storage[2562] = 0;
storage[2563] = 0;
storage[2564] = 0;
storage[2565] = 0;
storage[2566] = 0;
storage[2567] = 0;
storage[2568] = 0;
storage[2569] = 0;
storage[2570] = 0;
storage[2571] = 0;
storage[2572] = 0;
storage[2573] = 0;
storage[2574] = 0;
storage[2575] = 0;
storage[2576] = 0;
storage[2577] = 0;
storage[2578] = 0;
storage[2579] = 0;
storage[2580] = 0;
storage[2581] = 0;
storage[2582] = 0;
storage[2583] = 0;
storage[2584] = 0;
storage[2585] = 0;
storage[2586] = 0;
storage[2587] = 0;
storage[2588] = 0;
storage[2589] = 0;
storage[2590] = 0;
storage[2591] = 0;
storage[2592] = 0;
storage[2593] = 0;
storage[2594] = 0;
storage[2595] = 0;
storage[2596] = 0;
storage[2597] = 0;
storage[2598] = 0;
storage[2599] = 0;
storage[2600] = 0;
storage[2601] = 0;
storage[2602] = 0;
storage[2603] = 0;
storage[2604] = 0;
storage[2605] = 0;
storage[2606] = 0;
storage[2607] = 0;
storage[2608] = 0;
storage[2609] = 0;
storage[2610] = 0;
storage[2611] = 0;
storage[2612] = 0;
storage[2613] = 0;
storage[2614] = 0;
storage[2615] = 0;
storage[2616] = 0;
storage[2617] = 0;
storage[2618] = 0;
storage[2619] = 0;
storage[2620] = 0;
storage[2621] = 0;
storage[2622] = 0;
storage[2623] = 0;
storage[2624] = 0;
storage[2625] = 0;
storage[2626] = 0;
storage[2627] = 0;
storage[2628] = 0;
storage[2629] = 0;
storage[2630] = 0;
storage[2631] = 0;
storage[2632] = 0;
storage[2633] = 0;
storage[2634] = 0;
storage[2635] = 0;
storage[2636] = 0;
storage[2637] = 0;
storage[2638] = 0;
storage[2639] = 0;
storage[2640] = 0;
storage[2641] = 0;
storage[2642] = 0;
storage[2643] = 0;
storage[2644] = 0;
storage[2645] = 0;
storage[2646] = 0;
storage[2647] = 0;
storage[2648] = 0;
storage[2649] = 0;
storage[2650] = 0;
storage[2651] = 0;
storage[2652] = 0;
storage[2653] = 0;
storage[2654] = 0;
storage[2655] = 0;
storage[2656] = 0;
storage[2657] = 0;
storage[2658] = 0;
storage[2659] = 0;
storage[2660] = 0;
storage[2661] = 0;
storage[2662] = 0;
storage[2663] = 0;
storage[2664] = 0;
storage[2665] = 0;
storage[2666] = 0;
storage[2667] = 0;
storage[2668] = 0;
storage[2669] = 0;
storage[2670] = 0;
storage[2671] = 0;
storage[2672] = 0;
storage[2673] = 0;
storage[2674] = 0;
storage[2675] = 0;
storage[2676] = 0;
storage[2677] = 0;
storage[2678] = 0;
storage[2679] = 0;
storage[2680] = 0;
storage[2681] = 0;
storage[2682] = 0;
storage[2683] = 0;
storage[2684] = 0;
storage[2685] = 0;
storage[2686] = 0;
storage[2687] = 0;
storage[2688] = 0;
storage[2689] = 0;
storage[2690] = 0;
storage[2691] = 0;
storage[2692] = 0;
storage[2693] = 0;
storage[2694] = 0;
storage[2695] = 0;
storage[2696] = 0;
storage[2697] = 0;
storage[2698] = 0;
storage[2699] = 0;
storage[2700] = 0;
storage[2701] = 0;
storage[2702] = 0;
storage[2703] = 0;
storage[2704] = 0;
storage[2705] = 0;
storage[2706] = 0;
storage[2707] = 0;
storage[2708] = 0;
storage[2709] = 0;
storage[2710] = 0;
storage[2711] = 0;
storage[2712] = 0;
storage[2713] = 0;
storage[2714] = 0;
storage[2715] = 0;
storage[2716] = 0;
storage[2717] = 0;
storage[2718] = 0;
storage[2719] = 0;
storage[2720] = 0;
storage[2721] = 0;
storage[2722] = 0;
storage[2723] = 0;
storage[2724] = 0;
storage[2725] = 0;
storage[2726] = 0;
storage[2727] = 0;
storage[2728] = 0;
storage[2729] = 0;
storage[2730] = 0;
storage[2731] = 0;
storage[2732] = 0;
storage[2733] = 0;
storage[2734] = 0;
storage[2735] = 0;
storage[2736] = 0;
storage[2737] = 0;
storage[2738] = 0;
storage[2739] = 0;
storage[2740] = 0;
storage[2741] = 0;
storage[2742] = 0;
storage[2743] = 0;
storage[2744] = 0;
storage[2745] = 0;
storage[2746] = 0;
storage[2747] = 0;
storage[2748] = 0;
storage[2749] = 0;
storage[2750] = 0;
storage[2751] = 0;
storage[2752] = 0;
storage[2753] = 0;
storage[2754] = 0;
storage[2755] = 0;
storage[2756] = 0;
storage[2757] = 0;
storage[2758] = 0;
storage[2759] = 0;
storage[2760] = 0;
storage[2761] = 0;
storage[2762] = 0;
storage[2763] = 0;
storage[2764] = 0;
storage[2765] = 0;
storage[2766] = 0;
storage[2767] = 0;
storage[2768] = 0;
storage[2769] = 0;
storage[2770] = 0;
storage[2771] = 0;
storage[2772] = 0;
storage[2773] = 0;
storage[2774] = 0;
storage[2775] = 0;
storage[2776] = 0;
storage[2777] = 0;
storage[2778] = 0;
storage[2779] = 0;
storage[2780] = 0;
storage[2781] = 0;
storage[2782] = 0;
storage[2783] = 0;
storage[2784] = 0;
storage[2785] = 0;
storage[2786] = 0;
storage[2787] = 0;
storage[2788] = 0;
storage[2789] = 0;
storage[2790] = 0;
storage[2791] = 0;
storage[2792] = 0;
storage[2793] = 0;
storage[2794] = 0;
storage[2795] = 0;
storage[2796] = 0;
storage[2797] = 0;
storage[2798] = 0;
storage[2799] = 0;
storage[2800] = 0;
storage[2801] = 0;
storage[2802] = 0;
storage[2803] = 0;
storage[2804] = 0;
storage[2805] = 0;
storage[2806] = 0;
storage[2807] = 0;
storage[2808] = 0;
storage[2809] = 0;
storage[2810] = 0;
storage[2811] = 0;
storage[2812] = 0;
storage[2813] = 0;
storage[2814] = 0;
storage[2815] = 0;
storage[2816] = 0;
storage[2817] = 0;
storage[2818] = 0;
storage[2819] = 0;
storage[2820] = 0;
storage[2821] = 0;
storage[2822] = 0;
storage[2823] = 0;
storage[2824] = 0;
storage[2825] = 0;
storage[2826] = 0;
storage[2827] = 0;
storage[2828] = 0;
storage[2829] = 0;
storage[2830] = 0;
storage[2831] = 0;
storage[2832] = 0;
storage[2833] = 0;
storage[2834] = 0;
storage[2835] = 0;
storage[2836] = 0;
storage[2837] = 0;
storage[2838] = 0;
storage[2839] = 0;
storage[2840] = 0;
storage[2841] = 0;
storage[2842] = 0;
storage[2843] = 0;
storage[2844] = 0;
storage[2845] = 0;
storage[2846] = 0;
storage[2847] = 0;
storage[2848] = 0;
storage[2849] = 0;
storage[2850] = 0;
storage[2851] = 0;
storage[2852] = 0;
storage[2853] = 0;
storage[2854] = 0;
storage[2855] = 0;
storage[2856] = 0;
storage[2857] = 0;
storage[2858] = 0;
storage[2859] = 0;
storage[2860] = 0;
storage[2861] = 0;
storage[2862] = 0;
storage[2863] = 0;
storage[2864] = 0;
storage[2865] = 0;
storage[2866] = 0;
storage[2867] = 0;
storage[2868] = 0;
storage[2869] = 0;
storage[2870] = 0;
storage[2871] = 0;
storage[2872] = 0;
storage[2873] = 0;
storage[2874] = 0;
storage[2875] = 0;
storage[2876] = 0;
storage[2877] = 0;
storage[2878] = 0;
storage[2879] = 0;
storage[2880] = 0;
storage[2881] = 0;
storage[2882] = 0;
storage[2883] = 0;
storage[2884] = 0;
storage[2885] = 0;
storage[2886] = 0;
storage[2887] = 0;
storage[2888] = 0;
storage[2889] = 0;
storage[2890] = 0;
storage[2891] = 0;
storage[2892] = 0;
storage[2893] = 0;
storage[2894] = 0;
storage[2895] = 0;
storage[2896] = 0;
storage[2897] = 0;
storage[2898] = 0;
storage[2899] = 0;
storage[2900] = 0;
storage[2901] = 0;
storage[2902] = 0;
storage[2903] = 0;
storage[2904] = 0;
storage[2905] = 0;
storage[2906] = 0;
storage[2907] = 0;
storage[2908] = 0;
storage[2909] = 0;
storage[2910] = 0;
storage[2911] = 0;
storage[2912] = 0;
storage[2913] = 0;
storage[2914] = 0;
storage[2915] = 0;
storage[2916] = 0;
storage[2917] = 0;
storage[2918] = 0;
storage[2919] = 0;
storage[2920] = 0;
storage[2921] = 0;
storage[2922] = 0;
storage[2923] = 0;
storage[2924] = 0;
storage[2925] = 0;
storage[2926] = 0;
storage[2927] = 0;
storage[2928] = 0;
storage[2929] = 0;
storage[2930] = 0;
storage[2931] = 0;
storage[2932] = 0;
storage[2933] = 0;
storage[2934] = 0;
storage[2935] = 0;
storage[2936] = 0;
storage[2937] = 0;
storage[2938] = 0;
storage[2939] = 0;
storage[2940] = 0;
storage[2941] = 0;
storage[2942] = 0;
storage[2943] = 0;
storage[2944] = 0;
storage[2945] = 0;
storage[2946] = 0;
storage[2947] = 0;
storage[2948] = 0;
storage[2949] = 0;
storage[2950] = 0;
storage[2951] = 0;
storage[2952] = 0;
storage[2953] = 0;
storage[2954] = 0;
storage[2955] = 0;
storage[2956] = 0;
storage[2957] = 0;
storage[2958] = 0;
storage[2959] = 0;
storage[2960] = 0;
storage[2961] = 0;
storage[2962] = 0;
storage[2963] = 0;
storage[2964] = 0;
storage[2965] = 0;
storage[2966] = 0;
storage[2967] = 0;
storage[2968] = 0;
storage[2969] = 0;
storage[2970] = 0;
storage[2971] = 0;
storage[2972] = 0;
storage[2973] = 0;
storage[2974] = 0;
storage[2975] = 0;
storage[2976] = 0;
storage[2977] = 0;
storage[2978] = 0;
storage[2979] = 0;
storage[2980] = 0;
storage[2981] = 0;
storage[2982] = 0;
storage[2983] = 0;
storage[2984] = 0;
storage[2985] = 0;
storage[2986] = 0;
storage[2987] = 0;
storage[2988] = 0;
storage[2989] = 0;
storage[2990] = 0;
storage[2991] = 0;
storage[2992] = 0;
storage[2993] = 0;
storage[2994] = 0;
storage[2995] = 0;
storage[2996] = 0;
storage[2997] = 0;
storage[2998] = 0;
storage[2999] = 0;
storage[3000] = 0;
storage[3001] = 0;
storage[3002] = 0;
storage[3003] = 0;
storage[3004] = 0;
storage[3005] = 0;
storage[3006] = 0;
storage[3007] = 0;
storage[3008] = 0;
storage[3009] = 0;
storage[3010] = 0;
storage[3011] = 0;
storage[3012] = 0;
storage[3013] = 0;
storage[3014] = 0;
storage[3015] = 0;
storage[3016] = 0;
storage[3017] = 0;
storage[3018] = 0;
storage[3019] = 0;
storage[3020] = 0;
storage[3021] = 0;
storage[3022] = 0;
storage[3023] = 0;
storage[3024] = 0;
storage[3025] = 0;
storage[3026] = 0;
storage[3027] = 0;
storage[3028] = 0;
storage[3029] = 0;
storage[3030] = 0;
storage[3031] = 0;
storage[3032] = 0;
storage[3033] = 0;
storage[3034] = 0;
storage[3035] = 0;
storage[3036] = 0;
storage[3037] = 0;
storage[3038] = 0;
storage[3039] = 0;
storage[3040] = 0;
storage[3041] = 0;
storage[3042] = 0;
storage[3043] = 0;
storage[3044] = 0;
storage[3045] = 0;
storage[3046] = 0;
storage[3047] = 0;
storage[3048] = 0;
storage[3049] = 0;
storage[3050] = 0;
storage[3051] = 0;
storage[3052] = 0;
storage[3053] = 0;
storage[3054] = 0;
storage[3055] = 0;
storage[3056] = 0;
storage[3057] = 0;
storage[3058] = 0;
storage[3059] = 0;
storage[3060] = 0;
storage[3061] = 0;
storage[3062] = 0;
storage[3063] = 0;
storage[3064] = 0;
storage[3065] = 0;
storage[3066] = 0;
storage[3067] = 0;
storage[3068] = 0;
storage[3069] = 0;
storage[3070] = 0;
storage[3071] = 0;
storage[3072] = 0;
storage[3073] = 0;
storage[3074] = 0;
storage[3075] = 0;
storage[3076] = 0;
storage[3077] = 0;
storage[3078] = 0;
storage[3079] = 0;
storage[3080] = 0;
storage[3081] = 0;
storage[3082] = 0;
storage[3083] = 0;
storage[3084] = 0;
storage[3085] = 0;
storage[3086] = 0;
storage[3087] = 0;
storage[3088] = 0;
storage[3089] = 0;
storage[3090] = 0;
storage[3091] = 0;
storage[3092] = 0;
storage[3093] = 0;
storage[3094] = 0;
storage[3095] = 0;
storage[3096] = 0;
storage[3097] = 0;
storage[3098] = 0;
storage[3099] = 0;
storage[3100] = 0;
storage[3101] = 0;
storage[3102] = 0;
storage[3103] = 0;
storage[3104] = 0;
storage[3105] = 0;
storage[3106] = 0;
storage[3107] = 0;
storage[3108] = 0;
storage[3109] = 0;
storage[3110] = 0;
storage[3111] = 0;
storage[3112] = 0;
storage[3113] = 0;
storage[3114] = 0;
storage[3115] = 0;
storage[3116] = 0;
storage[3117] = 0;
storage[3118] = 0;
storage[3119] = 0;
storage[3120] = 0;
storage[3121] = 0;
storage[3122] = 0;
storage[3123] = 0;
storage[3124] = 0;
storage[3125] = 0;
storage[3126] = 0;
storage[3127] = 0;
storage[3128] = 0;
storage[3129] = 0;
storage[3130] = 0;
storage[3131] = 0;
storage[3132] = 0;
storage[3133] = 0;
storage[3134] = 0;
storage[3135] = 0;
storage[3136] = 0;
storage[3137] = 0;
storage[3138] = 0;
storage[3139] = 0;
storage[3140] = 0;
storage[3141] = 0;
storage[3142] = 0;
storage[3143] = 0;
storage[3144] = 0;
storage[3145] = 0;
storage[3146] = 0;
storage[3147] = 0;
storage[3148] = 0;
storage[3149] = 0;
storage[3150] = 0;
storage[3151] = 0;
storage[3152] = 0;
storage[3153] = 0;
storage[3154] = 0;
storage[3155] = 0;
storage[3156] = 0;
storage[3157] = 0;
storage[3158] = 0;
storage[3159] = 0;
storage[3160] = 0;
storage[3161] = 0;
storage[3162] = 0;
storage[3163] = 0;
storage[3164] = 0;
storage[3165] = 0;
storage[3166] = 0;
storage[3167] = 0;
storage[3168] = 0;
storage[3169] = 0;
storage[3170] = 0;
storage[3171] = 0;
storage[3172] = 0;
storage[3173] = 0;
storage[3174] = 0;
storage[3175] = 0;
storage[3176] = 0;
storage[3177] = 0;
storage[3178] = 0;
storage[3179] = 0;
storage[3180] = 0;
storage[3181] = 0;
storage[3182] = 0;
storage[3183] = 0;
storage[3184] = 0;
storage[3185] = 0;
storage[3186] = 0;
storage[3187] = 0;
storage[3188] = 0;
storage[3189] = 0;
storage[3190] = 0;
storage[3191] = 0;
storage[3192] = 0;
storage[3193] = 0;
storage[3194] = 0;
storage[3195] = 0;
storage[3196] = 0;
storage[3197] = 0;
storage[3198] = 0;
storage[3199] = 0;   
	end

	always @(posedge clk) begin
		if(we==1) begin
			storage[address_p+1] <= dp;
		end
	end
		
	always @(posedge clk) begin
		if(re==1) begin
			datata <= storage[address];
		end
    end
endmodule
