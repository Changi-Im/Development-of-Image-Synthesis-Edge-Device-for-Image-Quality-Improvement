module test();

  parameter SIZE=14;

  reg clk;
  reg GO;
  reg signed [SIZE-1:0] storage1 [0:3199]; 
  wire STOP;
  
  reg we_database;
  reg [SIZE-1:0] dp_database;
  reg [15:0] address_p_database;
  
  reg [13:0] x;
  
  wire signed [13:0] image_final;
  wire                  image_final_en;
  
  TOP TOP(
	.clk					(clk),
	.GO						(GO),
	.we_database			(we_database), 
	.dp_database			(dp_database), 
	.address_p_database		(address_p_database-1'b1),
	.STOP					(STOP),
	.image_final            (image_final),
	.image_final_en         (image_final_en)
  );
      
    initial begin
      clk                = 0;
      address_p_database = 0;
      x                  = 0;
      we_database        = 1;
      #200 GO            = 1;
    end
    
    always #1 clk = ~clk;
    
    always @(posedge clk) begin
        if(we_database) begin
            if(address_p_database<=3199) begin
                dp_database = storage1[address_p_database];
                address_p_database=address_p_database+1'b1;
            end else begin
                we_database=0;
            end 
        end
        
        if((x<=40*40*2)&&(GO)) begin
            x=x+1;
        end else begin
            GO=0;
        end
        
        if(STOP==1) begin
           $finish;
        end
        
        if(image_final_en == 1) begin   
            #32 $display("'0b%b',",image_final);
        end
     end
     
   initial begin
    // image 1
storage1[0] = 14'b000000000_0000;
storage1[1] = 14'b000000000_0000;
storage1[2] = 14'b000000000_0000;
storage1[3] = 14'b000000001_0000;
storage1[4] = 14'b000000000_0000;
storage1[5] = 14'b000000000_0000;
storage1[6] = 14'b000000000_0000;
storage1[7] = 14'b000000001_0000;
storage1[8] = 14'b000000000_0000;
storage1[9] = 14'b000000000_0000;
storage1[10] = 14'b000000000_0000;
storage1[11] = 14'b000000001_0000;
storage1[12] = 14'b000000001_0000;
storage1[13] = 14'b000000001_0000;
storage1[14] = 14'b000000001_0000;
storage1[15] = 14'b000000001_0000;
storage1[16] = 14'b000000001_0000;
storage1[17] = 14'b000000001_0000;
storage1[18] = 14'b000000001_0000;
storage1[19] = 14'b000000001_0000;
storage1[20] = 14'b000000000_0000;
storage1[21] = 14'b000000000_0000;
storage1[22] = 14'b000000000_0000;
storage1[23] = 14'b000000000_0000;
storage1[24] = 14'b000000000_0000;
storage1[25] = 14'b000000000_0000;
storage1[26] = 14'b000000111_0000;
storage1[27] = 14'b001011110_0000;
storage1[28] = 14'b000001001_0000;
storage1[29] = 14'b000000001_0000;
storage1[30] = 14'b000000000_0000;
storage1[31] = 14'b000000001_0000;
storage1[32] = 14'b000000000_0000;
storage1[33] = 14'b000000000_0000;
storage1[34] = 14'b000000000_0000;
storage1[35] = 14'b000000000_0000;
storage1[36] = 14'b000000000_0000;
storage1[37] = 14'b000000001_0000;
storage1[38] = 14'b000000000_0000;
storage1[39] = 14'b000000000_0000;
storage1[40] = 14'b000000000_0000;
storage1[41] = 14'b000000000_0000;
storage1[42] = 14'b000000000_0000;
storage1[43] = 14'b000000000_0000;
storage1[44] = 14'b000000000_0000;
storage1[45] = 14'b000000000_0000;
storage1[46] = 14'b000000000_0000;
storage1[47] = 14'b000000000_0000;
storage1[48] = 14'b000000000_0000;
storage1[49] = 14'b000000000_0000;
storage1[50] = 14'b000000000_0000;
storage1[51] = 14'b000000000_0000;
storage1[52] = 14'b000000000_0000;
storage1[53] = 14'b000000000_0000;
storage1[54] = 14'b000000000_0000;
storage1[55] = 14'b000000001_0000;
storage1[56] = 14'b000000000_0000;
storage1[57] = 14'b000000000_0000;
storage1[58] = 14'b000000001_0000;
storage1[59] = 14'b000000000_0000;
storage1[60] = 14'b000000000_0000;
storage1[61] = 14'b000000001_0000;
storage1[62] = 14'b000000000_0000;
storage1[63] = 14'b000000000_0000;
storage1[64] = 14'b000000000_0000;
storage1[65] = 14'b000000001_0000;
storage1[66] = 14'b000000000_0000;
storage1[67] = 14'b000000011_0000;
storage1[68] = 14'b000000001_0000;
storage1[69] = 14'b000000001_0000;
storage1[70] = 14'b000000000_0000;
storage1[71] = 14'b000000000_0000;
storage1[72] = 14'b000000000_0000;
storage1[73] = 14'b000000000_0000;
storage1[74] = 14'b000000000_0000;
storage1[75] = 14'b000000000_0000;
storage1[76] = 14'b000000000_0000;
storage1[77] = 14'b000000000_0000;
storage1[78] = 14'b000000000_0000;
storage1[79] = 14'b000000000_0000;
storage1[80] = 14'b000000001_0000;
storage1[81] = 14'b000000010_0000;
storage1[82] = 14'b000000001_0000;
storage1[83] = 14'b000000010_0000;
storage1[84] = 14'b000000010_0000;
storage1[85] = 14'b000000001_0000;
storage1[86] = 14'b000000010_0000;
storage1[87] = 14'b000000001_0000;
storage1[88] = 14'b000000010_0000;
storage1[89] = 14'b000000010_0000;
storage1[90] = 14'b000000010_0000;
storage1[91] = 14'b000000010_0000;
storage1[92] = 14'b000000011_0000;
storage1[93] = 14'b000000010_0000;
storage1[94] = 14'b000000011_0000;
storage1[95] = 14'b000000101_0000;
storage1[96] = 14'b000000010_0000;
storage1[97] = 14'b000000011_0000;
storage1[98] = 14'b000000010_0000;
storage1[99] = 14'b000000101_0000;
storage1[100] = 14'b000000010_0000;
storage1[101] = 14'b000000011_0000;
storage1[102] = 14'b000000011_0000;
storage1[103] = 14'b000000011_0000;
storage1[104] = 14'b000000011_0000;
storage1[105] = 14'b000000101_0000;
storage1[106] = 14'b000000010_0000;
storage1[107] = 14'b000000010_0000;
storage1[108] = 14'b000000011_0000;
storage1[109] = 14'b000000011_0000;
storage1[110] = 14'b000000010_0000;
storage1[111] = 14'b000000001_0000;
storage1[112] = 14'b000000000_0000;
storage1[113] = 14'b000000000_0000;
storage1[114] = 14'b000000000_0000;
storage1[115] = 14'b000000000_0000;
storage1[116] = 14'b000000000_0000;
storage1[117] = 14'b000000000_0000;
storage1[118] = 14'b000000000_0000;
storage1[119] = 14'b000000000_0000;
storage1[120] = 14'b000000010_0000;
storage1[121] = 14'b000000010_0000;
storage1[122] = 14'b000000001_0000;
storage1[123] = 14'b000000010_0000;
storage1[124] = 14'b000000011_0000;
storage1[125] = 14'b000000011_0000;
storage1[126] = 14'b000000010_0000;
storage1[127] = 14'b000000011_0000;
storage1[128] = 14'b000000010_0000;
storage1[129] = 14'b000000010_0000;
storage1[130] = 14'b000000010_0000;
storage1[131] = 14'b000000010_0000;
storage1[132] = 14'b000000011_0000;
storage1[133] = 14'b000000010_0000;
storage1[134] = 14'b000000011_0000;
storage1[135] = 14'b000000011_0000;
storage1[136] = 14'b000000011_0000;
storage1[137] = 14'b000000011_0000;
storage1[138] = 14'b000000011_0000;
storage1[139] = 14'b000000011_0000;
storage1[140] = 14'b000000010_0000;
storage1[141] = 14'b000000011_0000;
storage1[142] = 14'b000000101_0000;
storage1[143] = 14'b000000011_0000;
storage1[144] = 14'b000000010_0000;
storage1[145] = 14'b000000011_0000;
storage1[146] = 14'b000000010_0000;
storage1[147] = 14'b000000011_0000;
storage1[148] = 14'b000000101_0000;
storage1[149] = 14'b000000010_0000;
storage1[150] = 14'b000000010_0000;
storage1[151] = 14'b000000001_0000;
storage1[152] = 14'b000000000_0000;
storage1[153] = 14'b000000001_0000;
storage1[154] = 14'b000000001_0000;
storage1[155] = 14'b000000001_0000;
storage1[156] = 14'b000000000_0000;
storage1[157] = 14'b000000000_0000;
storage1[158] = 14'b000000000_0000;
storage1[159] = 14'b000000000_0000;
storage1[160] = 14'b000000010_0000;
storage1[161] = 14'b000000010_0000;
storage1[162] = 14'b000000010_0000;
storage1[163] = 14'b000000001_0000;
storage1[164] = 14'b000000010_0000;
storage1[165] = 14'b000000010_0000;
storage1[166] = 14'b000000010_0000;
storage1[167] = 14'b000000010_0000;
storage1[168] = 14'b000000010_0000;
storage1[169] = 14'b000000011_0000;
storage1[170] = 14'b000000011_0000;
storage1[171] = 14'b000000010_0000;
storage1[172] = 14'b000000101_0000;
storage1[173] = 14'b000000101_0000;
storage1[174] = 14'b000000011_0000;
storage1[175] = 14'b000000011_0000;
storage1[176] = 14'b000000010_0000;
storage1[177] = 14'b000000011_0000;
storage1[178] = 14'b000000011_0000;
storage1[179] = 14'b000000011_0000;
storage1[180] = 14'b000000101_0000;
storage1[181] = 14'b000000101_0000;
storage1[182] = 14'b000000101_0000;
storage1[183] = 14'b000000101_0000;
storage1[184] = 14'b000000101_0000;
storage1[185] = 14'b000000101_0000;
storage1[186] = 14'b000000101_0000;
storage1[187] = 14'b000000101_0000;
storage1[188] = 14'b000000011_0000;
storage1[189] = 14'b000000011_0000;
storage1[190] = 14'b000000001_0000;
storage1[191] = 14'b000000001_0000;
storage1[192] = 14'b000000001_0000;
storage1[193] = 14'b000000001_0000;
storage1[194] = 14'b000001110_0000;
storage1[195] = 14'b000000001_0000;
storage1[196] = 14'b000000001_0000;
storage1[197] = 14'b000000000_0000;
storage1[198] = 14'b000000000_0000;
storage1[199] = 14'b000000001_0000;
storage1[200] = 14'b000000010_0000;
storage1[201] = 14'b000000011_0000;
storage1[202] = 14'b000000011_0000;
storage1[203] = 14'b000000010_0000;
storage1[204] = 14'b000000001_0000;
storage1[205] = 14'b000000010_0000;
storage1[206] = 14'b000000010_0000;
storage1[207] = 14'b000000010_0000;
storage1[208] = 14'b000000010_0000;
storage1[209] = 14'b000000010_0000;
storage1[210] = 14'b000000010_0000;
storage1[211] = 14'b000000010_0000;
storage1[212] = 14'b000000101_0000;
storage1[213] = 14'b000000101_0000;
storage1[214] = 14'b000000011_0000;
storage1[215] = 14'b000000011_0000;
storage1[216] = 14'b000000011_0000;
storage1[217] = 14'b000000011_0000;
storage1[218] = 14'b000000010_0000;
storage1[219] = 14'b000000011_0000;
storage1[220] = 14'b000000101_0000;
storage1[221] = 14'b000000101_0000;
storage1[222] = 14'b000000101_0000;
storage1[223] = 14'b000000011_0000;
storage1[224] = 14'b000000011_0000;
storage1[225] = 14'b000000010_0000;
storage1[226] = 14'b000000101_0000;
storage1[227] = 14'b000000101_0000;
storage1[228] = 14'b000000011_0000;
storage1[229] = 14'b000000101_0000;
storage1[230] = 14'b000000001_0000;
storage1[231] = 14'b000000001_0000;
storage1[232] = 14'b000000001_0000;
storage1[233] = 14'b000001110_0000;
storage1[234] = 14'b000111110_0000;
storage1[235] = 14'b000000001_0000;
storage1[236] = 14'b000000001_0000;
storage1[237] = 14'b000000000_0000;
storage1[238] = 14'b000000001_0000;
storage1[239] = 14'b000000000_0000;
storage1[240] = 14'b000000001_0000;
storage1[241] = 14'b000000011_0000;
storage1[242] = 14'b000000011_0000;
storage1[243] = 14'b000000010_0000;
storage1[244] = 14'b000000001_0000;
storage1[245] = 14'b000000001_0000;
storage1[246] = 14'b000000001_0000;
storage1[247] = 14'b000000011_0000;
storage1[248] = 14'b000000011_0000;
storage1[249] = 14'b000000001_0000;
storage1[250] = 14'b000000001_0000;
storage1[251] = 14'b000000001_0000;
storage1[252] = 14'b000000011_0000;
storage1[253] = 14'b000000011_0000;
storage1[254] = 14'b000000010_0000;
storage1[255] = 14'b000000010_0000;
storage1[256] = 14'b000000001_0000;
storage1[257] = 14'b000000010_0000;
storage1[258] = 14'b000000001_0000;
storage1[259] = 14'b000000010_0000;
storage1[260] = 14'b000000011_0000;
storage1[261] = 14'b000000101_0000;
storage1[262] = 14'b000000010_0000;
storage1[263] = 14'b000000001_0000;
storage1[264] = 14'b000000000_0000;
storage1[265] = 14'b000000001_0000;
storage1[266] = 14'b000000010_0000;
storage1[267] = 14'b000000011_0000;
storage1[268] = 14'b000000101_0000;
storage1[269] = 14'b000000011_0000;
storage1[270] = 14'b000000001_0000;
storage1[271] = 14'b000000001_0000;
storage1[272] = 14'b000000010_0000;
storage1[273] = 14'b000000010_0000;
storage1[274] = 14'b000010010_0000;
storage1[275] = 14'b000000001_0000;
storage1[276] = 14'b000000001_0000;
storage1[277] = 14'b000000000_0000;
storage1[278] = 14'b000000000_0000;
storage1[279] = 14'b000000000_0000;
storage1[280] = 14'b000000001_0000;
storage1[281] = 14'b000000010_0000;
storage1[282] = 14'b000000011_0000;
storage1[283] = 14'b000000011_0000;
storage1[284] = 14'b000000110_0000;
storage1[285] = 14'b000101110_0000;
storage1[286] = 14'b000000110_0000;
storage1[287] = 14'b000000101_0000;
storage1[288] = 14'b000000011_0000;
storage1[289] = 14'b000000001_0000;
storage1[290] = 14'b000000111_0000;
storage1[291] = 14'b000010000_0000;
storage1[292] = 14'b000000010_0000;
storage1[293] = 14'b000000101_0000;
storage1[294] = 14'b000000101_0000;
storage1[295] = 14'b000000010_0000;
storage1[296] = 14'b000000010_0000;
storage1[297] = 14'b000101011_0000;
storage1[298] = 14'b000010001_0000;
storage1[299] = 14'b000000010_0000;
storage1[300] = 14'b000000101_0000;
storage1[301] = 14'b000000101_0000;
storage1[302] = 14'b000000010_0000;
storage1[303] = 14'b000000000_0000;
storage1[304] = 14'b000000000_0000;
storage1[305] = 14'b000000001_0000;
storage1[306] = 14'b000000010_0000;
storage1[307] = 14'b000000011_0000;
storage1[308] = 14'b000000101_0000;
storage1[309] = 14'b000000011_0000;
storage1[310] = 14'b000000001_0000;
storage1[311] = 14'b000000001_0000;
storage1[312] = 14'b000000001_0000;
storage1[313] = 14'b000000001_0000;
storage1[314] = 14'b000000000_0000;
storage1[315] = 14'b000000000_0000;
storage1[316] = 14'b000000000_0000;
storage1[317] = 14'b000000000_0000;
storage1[318] = 14'b000000000_0000;
storage1[319] = 14'b000000001_0000;
storage1[320] = 14'b000000001_0000;
storage1[321] = 14'b000000011_0000;
storage1[322] = 14'b000000010_0000;
storage1[323] = 14'b000000011_0000;
storage1[324] = 14'b000000101_0000;
storage1[325] = 14'b000011101_0000;
storage1[326] = 14'b000000101_0000;
storage1[327] = 14'b000000101_0000;
storage1[328] = 14'b000000011_0000;
storage1[329] = 14'b000000010_0000;
storage1[330] = 14'b000001001_0000;
storage1[331] = 14'b000001001_0000;
storage1[332] = 14'b000000010_0000;
storage1[333] = 14'b000000011_0000;
storage1[334] = 14'b000000011_0000;
storage1[335] = 14'b000000010_0000;
storage1[336] = 14'b000000001_0000;
storage1[337] = 14'b000011000_0000;
storage1[338] = 14'b000001001_0000;
storage1[339] = 14'b000000011_0000;
storage1[340] = 14'b000000011_0000;
storage1[341] = 14'b000000011_0000;
storage1[342] = 14'b000000001_0000;
storage1[343] = 14'b000000000_0000;
storage1[344] = 14'b000000000_0000;
storage1[345] = 14'b000000001_0000;
storage1[346] = 14'b000000010_0000;
storage1[347] = 14'b000000101_0000;
storage1[348] = 14'b000000011_0000;
storage1[349] = 14'b000000101_0000;
storage1[350] = 14'b000000001_0000;
storage1[351] = 14'b000000001_0000;
storage1[352] = 14'b000000001_0000;
storage1[353] = 14'b000000001_0000;
storage1[354] = 14'b000000001_0000;
storage1[355] = 14'b000000001_0000;
storage1[356] = 14'b000000001_0000;
storage1[357] = 14'b000000001_0000;
storage1[358] = 14'b000000000_0000;
storage1[359] = 14'b000000000_0000;
storage1[360] = 14'b000000000_0000;
storage1[361] = 14'b000000010_0000;
storage1[362] = 14'b000000010_0000;
storage1[363] = 14'b000000010_0000;
storage1[364] = 14'b000000001_0000;
storage1[365] = 14'b000000001_0000;
storage1[366] = 14'b000000001_0000;
storage1[367] = 14'b000000101_0000;
storage1[368] = 14'b000000011_0000;
storage1[369] = 14'b000000001_0000;
storage1[370] = 14'b000000001_0000;
storage1[371] = 14'b000000001_0000;
storage1[372] = 14'b000000010_0000;
storage1[373] = 14'b000000011_0000;
storage1[374] = 14'b000000101_0000;
storage1[375] = 14'b000000001_0000;
storage1[376] = 14'b000000001_0000;
storage1[377] = 14'b000000001_0000;
storage1[378] = 14'b000000001_0000;
storage1[379] = 14'b000000010_0000;
storage1[380] = 14'b000000101_0000;
storage1[381] = 14'b000000011_0000;
storage1[382] = 14'b000000010_0000;
storage1[383] = 14'b000000000_0000;
storage1[384] = 14'b000000000_0000;
storage1[385] = 14'b000000000_0000;
storage1[386] = 14'b000000010_0000;
storage1[387] = 14'b000000011_0000;
storage1[388] = 14'b000000101_0000;
storage1[389] = 14'b000000101_0000;
storage1[390] = 14'b000000010_0000;
storage1[391] = 14'b000000001_0000;
storage1[392] = 14'b000000001_0000;
storage1[393] = 14'b000000001_0000;
storage1[394] = 14'b000000001_0000;
storage1[395] = 14'b000000001_0000;
storage1[396] = 14'b000000001_0000;
storage1[397] = 14'b000000001_0000;
storage1[398] = 14'b000000000_0000;
storage1[399] = 14'b000000001_0000;
storage1[400] = 14'b000000001_0000;
storage1[401] = 14'b000000010_0000;
storage1[402] = 14'b000000011_0000;
storage1[403] = 14'b000000010_0000;
storage1[404] = 14'b000000001_0000;
storage1[405] = 14'b000000001_0000;
storage1[406] = 14'b000000001_0000;
storage1[407] = 14'b000000011_0000;
storage1[408] = 14'b000000011_0000;
storage1[409] = 14'b000000000_0000;
storage1[410] = 14'b000000001_0000;
storage1[411] = 14'b000000001_0000;
storage1[412] = 14'b000000011_0000;
storage1[413] = 14'b000000101_0000;
storage1[414] = 14'b000000101_0000;
storage1[415] = 14'b000000001_0000;
storage1[416] = 14'b000000001_0000;
storage1[417] = 14'b000000001_0000;
storage1[418] = 14'b000000001_0000;
storage1[419] = 14'b000000010_0000;
storage1[420] = 14'b000000011_0000;
storage1[421] = 14'b000000011_0000;
storage1[422] = 14'b000000001_0000;
storage1[423] = 14'b000000001_0000;
storage1[424] = 14'b000000010_0000;
storage1[425] = 14'b000000000_0000;
storage1[426] = 14'b000000010_0000;
storage1[427] = 14'b000000101_0000;
storage1[428] = 14'b000000101_0000;
storage1[429] = 14'b000000010_0000;
storage1[430] = 14'b000000001_0000;
storage1[431] = 14'b000000001_0000;
storage1[432] = 14'b000000001_0000;
storage1[433] = 14'b000000001_0000;
storage1[434] = 14'b000000001_0000;
storage1[435] = 14'b000000001_0000;
storage1[436] = 14'b000000001_0000;
storage1[437] = 14'b000000001_0000;
storage1[438] = 14'b000000000_0000;
storage1[439] = 14'b000000000_0000;
storage1[440] = 14'b000000000_0000;
storage1[441] = 14'b000000011_0000;
storage1[442] = 14'b000000010_0000;
storage1[443] = 14'b000000010_0000;
storage1[444] = 14'b000000010_0000;
storage1[445] = 14'b000001011_0000;
storage1[446] = 14'b000000111_0000;
storage1[447] = 14'b000000101_0000;
storage1[448] = 14'b000000010_0000;
storage1[449] = 14'b000000001_0000;
storage1[450] = 14'b000000101_0000;
storage1[451] = 14'b000000101_0000;
storage1[452] = 14'b000000011_0000;
storage1[453] = 14'b000000101_0000;
storage1[454] = 14'b000000101_0000;
storage1[455] = 14'b000000111_0000;
storage1[456] = 14'b000001100_0000;
storage1[457] = 14'b000001000_0000;
storage1[458] = 14'b000001010_0000;
storage1[459] = 14'b000000101_0000;
storage1[460] = 14'b000000101_0000;
storage1[461] = 14'b000000101_0000;
storage1[462] = 14'b000000010_0000;
storage1[463] = 14'b000001111_0000;
storage1[464] = 14'b000110011_0000;
storage1[465] = 14'b000010010_0000;
storage1[466] = 14'b000000011_0000;
storage1[467] = 14'b000000101_0000;
storage1[468] = 14'b000000101_0000;
storage1[469] = 14'b000000011_0000;
storage1[470] = 14'b000000001_0000;
storage1[471] = 14'b000000001_0000;
storage1[472] = 14'b000000001_0000;
storage1[473] = 14'b000000001_0000;
storage1[474] = 14'b000000000_0000;
storage1[475] = 14'b000000000_0000;
storage1[476] = 14'b000000001_0000;
storage1[477] = 14'b000000001_0000;
storage1[478] = 14'b000000000_0000;
storage1[479] = 14'b000000000_0000;
storage1[480] = 14'b000000001_0000;
storage1[481] = 14'b000000011_0000;
storage1[482] = 14'b000000011_0000;
storage1[483] = 14'b000000010_0000;
storage1[484] = 14'b000000001_0000;
storage1[485] = 14'b000001111_0000;
storage1[486] = 14'b000001100_0000;
storage1[487] = 14'b000000101_0000;
storage1[488] = 14'b000000010_0000;
storage1[489] = 14'b000000010_0000;
storage1[490] = 14'b000110010_0000;
storage1[491] = 14'b000100010_0000;
storage1[492] = 14'b000000101_0000;
storage1[493] = 14'b000000010_0000;
storage1[494] = 14'b000000101_0000;
storage1[495] = 14'b000001011_0000;
storage1[496] = 14'b000100100_0000;
storage1[497] = 14'b000010010_0000;
storage1[498] = 14'b000100100_0000;
storage1[499] = 14'b000000101_0000;
storage1[500] = 14'b000000101_0000;
storage1[501] = 14'b000000101_0000;
storage1[502] = 14'b000000010_0000;
storage1[503] = 14'b000111010_0000;
storage1[504] = 14'b001101001_0000;
storage1[505] = 14'b000100110_0000;
storage1[506] = 14'b000000101_0000;
storage1[507] = 14'b000000101_0000;
storage1[508] = 14'b000000101_0000;
storage1[509] = 14'b000000011_0000;
storage1[510] = 14'b000000001_0000;
storage1[511] = 14'b000000001_0000;
storage1[512] = 14'b000000001_0000;
storage1[513] = 14'b000000000_0000;
storage1[514] = 14'b000000000_0000;
storage1[515] = 14'b000000000_0000;
storage1[516] = 14'b000000001_0000;
storage1[517] = 14'b000000000_0000;
storage1[518] = 14'b000000000_0000;
storage1[519] = 14'b000000000_0000;
storage1[520] = 14'b000000010_0000;
storage1[521] = 14'b000000011_0000;
storage1[522] = 14'b000000011_0000;
storage1[523] = 14'b000000010_0000;
storage1[524] = 14'b000000010_0000;
storage1[525] = 14'b000000101_0000;
storage1[526] = 14'b000000101_0000;
storage1[527] = 14'b000000010_0000;
storage1[528] = 14'b000000101_0000;
storage1[529] = 14'b000000010_0000;
storage1[530] = 14'b000001011_0000;
storage1[531] = 14'b000001001_0000;
storage1[532] = 14'b000000011_0000;
storage1[533] = 14'b000000101_0000;
storage1[534] = 14'b000000101_0000;
storage1[535] = 14'b000000110_0000;
storage1[536] = 14'b000001010_0000;
storage1[537] = 14'b000000101_0000;
storage1[538] = 14'b000011111_0000;
storage1[539] = 14'b000000011_0000;
storage1[540] = 14'b000000010_0000;
storage1[541] = 14'b000000101_0000;
storage1[542] = 14'b000000010_0000;
storage1[543] = 14'b000000101_0000;
storage1[544] = 14'b000001011_0000;
storage1[545] = 14'b000001001_0000;
storage1[546] = 14'b000000101_0000;
storage1[547] = 14'b000000101_0000;
storage1[548] = 14'b000000101_0000;
storage1[549] = 14'b000000011_0000;
storage1[550] = 14'b000000001_0000;
storage1[551] = 14'b000000000_0000;
storage1[552] = 14'b000000001_0000;
storage1[553] = 14'b000000000_0000;
storage1[554] = 14'b000000000_0000;
storage1[555] = 14'b000000000_0000;
storage1[556] = 14'b000000000_0000;
storage1[557] = 14'b000000000_0000;
storage1[558] = 14'b000000000_0000;
storage1[559] = 14'b000000000_0000;
storage1[560] = 14'b000000010_0000;
storage1[561] = 14'b000000010_0000;
storage1[562] = 14'b000000011_0000;
storage1[563] = 14'b000000010_0000;
storage1[564] = 14'b000000101_0000;
storage1[565] = 14'b000000101_0000;
storage1[566] = 14'b000000010_0000;
storage1[567] = 14'b000000101_0000;
storage1[568] = 14'b000000101_0000;
storage1[569] = 14'b000000011_0000;
storage1[570] = 14'b000000101_0000;
storage1[571] = 14'b000000101_0000;
storage1[572] = 14'b000000101_0000;
storage1[573] = 14'b000000011_0000;
storage1[574] = 14'b000000101_0000;
storage1[575] = 14'b000000101_0000;
storage1[576] = 14'b000000010_0000;
storage1[577] = 14'b000000101_0000;
storage1[578] = 14'b000000101_0000;
storage1[579] = 14'b000000101_0000;
storage1[580] = 14'b000000101_0000;
storage1[581] = 14'b000000011_0000;
storage1[582] = 14'b000000011_0000;
storage1[583] = 14'b000000101_0000;
storage1[584] = 14'b000000101_0000;
storage1[585] = 14'b000000101_0000;
storage1[586] = 14'b000000011_0000;
storage1[587] = 14'b000000010_0000;
storage1[588] = 14'b000000011_0000;
storage1[589] = 14'b000000101_0000;
storage1[590] = 14'b000000000_0000;
storage1[591] = 14'b000000001_0000;
storage1[592] = 14'b000000001_0000;
storage1[593] = 14'b000000001_0000;
storage1[594] = 14'b000000000_0000;
storage1[595] = 14'b000000000_0000;
storage1[596] = 14'b000000000_0000;
storage1[597] = 14'b000000000_0000;
storage1[598] = 14'b000000000_0000;
storage1[599] = 14'b000000000_0000;
storage1[600] = 14'b000000010_0000;
storage1[601] = 14'b000000010_0000;
storage1[602] = 14'b000000010_0000;
storage1[603] = 14'b000000010_0000;
storage1[604] = 14'b000000010_0000;
storage1[605] = 14'b000000010_0000;
storage1[606] = 14'b000000001_0000;
storage1[607] = 14'b000000101_0000;
storage1[608] = 14'b000000011_0000;
storage1[609] = 14'b000000010_0000;
storage1[610] = 14'b000000010_0000;
storage1[611] = 14'b000000010_0000;
storage1[612] = 14'b000000011_0000;
storage1[613] = 14'b000000101_0000;
storage1[614] = 14'b000000101_0000;
storage1[615] = 14'b000000010_0000;
storage1[616] = 14'b000000101_0000;
storage1[617] = 14'b000000011_0000;
storage1[618] = 14'b000000011_0000;
storage1[619] = 14'b000000101_0000;
storage1[620] = 14'b000000101_0000;
storage1[621] = 14'b000000110_0000;
storage1[622] = 14'b000000010_0000;
storage1[623] = 14'b000000010_0000;
storage1[624] = 14'b000000011_0000;
storage1[625] = 14'b000000010_0000;
storage1[626] = 14'b000000011_0000;
storage1[627] = 14'b000000101_0000;
storage1[628] = 14'b000000101_0000;
storage1[629] = 14'b000000011_0000;
storage1[630] = 14'b000000001_0000;
storage1[631] = 14'b000000000_0000;
storage1[632] = 14'b000000001_0000;
storage1[633] = 14'b000000001_0000;
storage1[634] = 14'b000000000_0000;
storage1[635] = 14'b000000001_0000;
storage1[636] = 14'b000000000_0000;
storage1[637] = 14'b000000000_0000;
storage1[638] = 14'b000000000_0000;
storage1[639] = 14'b000000000_0000;
storage1[640] = 14'b000000010_0000;
storage1[641] = 14'b000000011_0000;
storage1[642] = 14'b000000010_0000;
storage1[643] = 14'b000000010_0000;
storage1[644] = 14'b000000000_0000;
storage1[645] = 14'b000000000_0000;
storage1[646] = 14'b000000010_0000;
storage1[647] = 14'b000000011_0000;
storage1[648] = 14'b000000101_0000;
storage1[649] = 14'b000000001_0000;
storage1[650] = 14'b000000001_0000;
storage1[651] = 14'b000000001_0000;
storage1[652] = 14'b000000101_0000;
storage1[653] = 14'b000000101_0000;
storage1[654] = 14'b000000101_0000;
storage1[655] = 14'b000000001_0000;
storage1[656] = 14'b000000000_0000;
storage1[657] = 14'b000000001_0000;
storage1[658] = 14'b000000001_0000;
storage1[659] = 14'b000000101_0000;
storage1[660] = 14'b000000101_0000;
storage1[661] = 14'b000000101_0000;
storage1[662] = 14'b000000001_0000;
storage1[663] = 14'b000000001_0000;
storage1[664] = 14'b000000000_0000;
storage1[665] = 14'b000000001_0000;
storage1[666] = 14'b000000101_0000;
storage1[667] = 14'b000000101_0000;
storage1[668] = 14'b000000101_0000;
storage1[669] = 14'b000000010_0000;
storage1[670] = 14'b000000001_0000;
storage1[671] = 14'b000000001_0000;
storage1[672] = 14'b000000001_0000;
storage1[673] = 14'b000000001_0000;
storage1[674] = 14'b000000000_0000;
storage1[675] = 14'b000000000_0000;
storage1[676] = 14'b000000001_0000;
storage1[677] = 14'b000000000_0000;
storage1[678] = 14'b000000000_0000;
storage1[679] = 14'b000000000_0000;
storage1[680] = 14'b000000010_0000;
storage1[681] = 14'b000000011_0000;
storage1[682] = 14'b000000101_0000;
storage1[683] = 14'b000000010_0000;
storage1[684] = 14'b000000000_0000;
storage1[685] = 14'b000000000_0000;
storage1[686] = 14'b000000010_0000;
storage1[687] = 14'b000000011_0000;
storage1[688] = 14'b000000011_0000;
storage1[689] = 14'b000000001_0000;
storage1[690] = 14'b000000001_0000;
storage1[691] = 14'b000000001_0000;
storage1[692] = 14'b000000101_0000;
storage1[693] = 14'b000000101_0000;
storage1[694] = 14'b000000101_0000;
storage1[695] = 14'b000000010_0000;
storage1[696] = 14'b000000010_0000;
storage1[697] = 14'b000000001_0000;
storage1[698] = 14'b000000001_0000;
storage1[699] = 14'b000000101_0000;
storage1[700] = 14'b000000101_0000;
storage1[701] = 14'b000000101_0000;
storage1[702] = 14'b000000001_0000;
storage1[703] = 14'b000000001_0000;
storage1[704] = 14'b000000001_0000;
storage1[705] = 14'b000000001_0000;
storage1[706] = 14'b000000101_0000;
storage1[707] = 14'b000000101_0000;
storage1[708] = 14'b000000101_0000;
storage1[709] = 14'b000000010_0000;
storage1[710] = 14'b000000001_0000;
storage1[711] = 14'b000000001_0000;
storage1[712] = 14'b000000001_0000;
storage1[713] = 14'b000000001_0000;
storage1[714] = 14'b000000001_0000;
storage1[715] = 14'b000000001_0000;
storage1[716] = 14'b000000001_0000;
storage1[717] = 14'b000000001_0000;
storage1[718] = 14'b000000000_0000;
storage1[719] = 14'b000000000_0000;
storage1[720] = 14'b000000010_0000;
storage1[721] = 14'b000000011_0000;
storage1[722] = 14'b000000010_0000;
storage1[723] = 14'b000000011_0000;
storage1[724] = 14'b000000011_0000;
storage1[725] = 14'b000000101_0000;
storage1[726] = 14'b000000011_0000;
storage1[727] = 14'b000000101_0000;
storage1[728] = 14'b000000011_0000;
storage1[729] = 14'b000000101_0000;
storage1[730] = 14'b000000101_0000;
storage1[731] = 14'b000000101_0000;
storage1[732] = 14'b000000101_0000;
storage1[733] = 14'b000000101_0000;
storage1[734] = 14'b000000101_0000;
storage1[735] = 14'b000000101_0000;
storage1[736] = 14'b000000101_0000;
storage1[737] = 14'b000000101_0000;
storage1[738] = 14'b000000101_0000;
storage1[739] = 14'b000000101_0000;
storage1[740] = 14'b000000101_0000;
storage1[741] = 14'b000000110_0000;
storage1[742] = 14'b000000101_0000;
storage1[743] = 14'b000000101_0000;
storage1[744] = 14'b000000101_0000;
storage1[745] = 14'b000000101_0000;
storage1[746] = 14'b000000101_0000;
storage1[747] = 14'b000000101_0000;
storage1[748] = 14'b000000101_0000;
storage1[749] = 14'b000000010_0000;
storage1[750] = 14'b000000001_0000;
storage1[751] = 14'b000000000_0000;
storage1[752] = 14'b000000001_0000;
storage1[753] = 14'b000000001_0000;
storage1[754] = 14'b000000001_0000;
storage1[755] = 14'b000000001_0000;
storage1[756] = 14'b000000001_0000;
storage1[757] = 14'b000000000_0000;
storage1[758] = 14'b000000000_0000;
storage1[759] = 14'b000000000_0000;
storage1[760] = 14'b000000011_0000;
storage1[761] = 14'b000000101_0000;
storage1[762] = 14'b000000011_0000;
storage1[763] = 14'b000000011_0000;
storage1[764] = 14'b000000101_0000;
storage1[765] = 14'b000000011_0000;
storage1[766] = 14'b000000010_0000;
storage1[767] = 14'b000000101_0000;
storage1[768] = 14'b000000011_0000;
storage1[769] = 14'b000000101_0000;
storage1[770] = 14'b000000101_0000;
storage1[771] = 14'b000000011_0000;
storage1[772] = 14'b000000101_0000;
storage1[773] = 14'b000000101_0000;
storage1[774] = 14'b000000101_0000;
storage1[775] = 14'b000000101_0000;
storage1[776] = 14'b000000101_0000;
storage1[777] = 14'b000000101_0000;
storage1[778] = 14'b000000110_0000;
storage1[779] = 14'b000000101_0000;
storage1[780] = 14'b000000101_0000;
storage1[781] = 14'b000000111_0000;
storage1[782] = 14'b000000011_0000;
storage1[783] = 14'b000000101_0000;
storage1[784] = 14'b000000110_0000;
storage1[785] = 14'b000000011_0000;
storage1[786] = 14'b000000101_0000;
storage1[787] = 14'b000000101_0000;
storage1[788] = 14'b000000101_0000;
storage1[789] = 14'b000000010_0000;
storage1[790] = 14'b000000010_0000;
storage1[791] = 14'b000000001_0000;
storage1[792] = 14'b000000001_0000;
storage1[793] = 14'b000000001_0000;
storage1[794] = 14'b000000001_0000;
storage1[795] = 14'b000000001_0000;
storage1[796] = 14'b000000001_0000;
storage1[797] = 14'b000000000_0000;
storage1[798] = 14'b000000000_0000;
storage1[799] = 14'b000000000_0000;
storage1[800] = 14'b000000010_0000;
storage1[801] = 14'b000000010_0000;
storage1[802] = 14'b000000011_0000;
storage1[803] = 14'b000000010_0000;
storage1[804] = 14'b000000001_0000;
storage1[805] = 14'b000000000_0000;
storage1[806] = 14'b000000010_0000;
storage1[807] = 14'b000000011_0000;
storage1[808] = 14'b000000011_0000;
storage1[809] = 14'b000001010_0000;
storage1[810] = 14'b000001111_0000;
storage1[811] = 14'b000001011_0000;
storage1[812] = 14'b000000101_0000;
storage1[813] = 14'b000000101_0000;
storage1[814] = 14'b000000011_0000;
storage1[815] = 14'b000000101_0000;
storage1[816] = 14'b000000110_0000;
storage1[817] = 14'b000001111_0000;
storage1[818] = 14'b000001001_0000;
storage1[819] = 14'b000000101_0000;
storage1[820] = 14'b000000101_0000;
storage1[821] = 14'b000000101_0000;
storage1[822] = 14'b000000001_0000;
storage1[823] = 14'b000000001_0000;
storage1[824] = 14'b000000001_0000;
storage1[825] = 14'b000000001_0000;
storage1[826] = 14'b000000011_0000;
storage1[827] = 14'b000000011_0000;
storage1[828] = 14'b000000101_0000;
storage1[829] = 14'b000000010_0000;
storage1[830] = 14'b000000010_0000;
storage1[831] = 14'b000000001_0000;
storage1[832] = 14'b000000001_0000;
storage1[833] = 14'b000000001_0000;
storage1[834] = 14'b000000001_0000;
storage1[835] = 14'b000000000_0000;
storage1[836] = 14'b000000001_0000;
storage1[837] = 14'b000000001_0000;
storage1[838] = 14'b000000001_0000;
storage1[839] = 14'b000000001_0000;
storage1[840] = 14'b000000010_0000;
storage1[841] = 14'b000000011_0000;
storage1[842] = 14'b000000101_0000;
storage1[843] = 14'b000000010_0000;
storage1[844] = 14'b000000000_0000;
storage1[845] = 14'b000000000_0000;
storage1[846] = 14'b000000010_0000;
storage1[847] = 14'b000000011_0000;
storage1[848] = 14'b000000101_0000;
storage1[849] = 14'b000010101_0000;
storage1[850] = 14'b000010101_0000;
storage1[851] = 14'b000001010_0000;
storage1[852] = 14'b000000101_0000;
storage1[853] = 14'b000000101_0000;
storage1[854] = 14'b000000101_0000;
storage1[855] = 14'b000000110_0000;
storage1[856] = 14'b000000111_0000;
storage1[857] = 14'b000001001_0000;
storage1[858] = 14'b000001100_0000;
storage1[859] = 14'b000000101_0000;
storage1[860] = 14'b000000101_0000;
storage1[861] = 14'b000000101_0000;
storage1[862] = 14'b000000000_0000;
storage1[863] = 14'b000000001_0000;
storage1[864] = 14'b000000001_0000;
storage1[865] = 14'b000000001_0000;
storage1[866] = 14'b000000101_0000;
storage1[867] = 14'b000000101_0000;
storage1[868] = 14'b000000110_0000;
storage1[869] = 14'b000000010_0000;
storage1[870] = 14'b000000001_0000;
storage1[871] = 14'b000000001_0000;
storage1[872] = 14'b000000001_0000;
storage1[873] = 14'b000000000_0000;
storage1[874] = 14'b000000001_0000;
storage1[875] = 14'b000000000_0000;
storage1[876] = 14'b000000001_0000;
storage1[877] = 14'b000000001_0000;
storage1[878] = 14'b000000001_0000;
storage1[879] = 14'b000000000_0000;
storage1[880] = 14'b000000010_0000;
storage1[881] = 14'b000000011_0000;
storage1[882] = 14'b000000011_0000;
storage1[883] = 14'b000000010_0000;
storage1[884] = 14'b000000010_0000;
storage1[885] = 14'b000000010_0000;
storage1[886] = 14'b000000101_0000;
storage1[887] = 14'b000000101_0000;
storage1[888] = 14'b000000011_0000;
storage1[889] = 14'b000000101_0000;
storage1[890] = 14'b000000101_0000;
storage1[891] = 14'b000000101_0000;
storage1[892] = 14'b000000101_0000;
storage1[893] = 14'b000000101_0000;
storage1[894] = 14'b000000101_0000;
storage1[895] = 14'b000000101_0000;
storage1[896] = 14'b000000101_0000;
storage1[897] = 14'b000000010_0000;
storage1[898] = 14'b000000101_0000;
storage1[899] = 14'b000000101_0000;
storage1[900] = 14'b000000101_0000;
storage1[901] = 14'b000000101_0000;
storage1[902] = 14'b000000011_0000;
storage1[903] = 14'b000000011_0000;
storage1[904] = 14'b000000011_0000;
storage1[905] = 14'b000000011_0000;
storage1[906] = 14'b000000101_0000;
storage1[907] = 14'b000000101_0000;
storage1[908] = 14'b000000101_0000;
storage1[909] = 14'b000000010_0000;
storage1[910] = 14'b000000001_0000;
storage1[911] = 14'b000000001_0000;
storage1[912] = 14'b000000001_0000;
storage1[913] = 14'b000000000_0000;
storage1[914] = 14'b000000000_0000;
storage1[915] = 14'b000000001_0000;
storage1[916] = 14'b000000001_0000;
storage1[917] = 14'b000000001_0000;
storage1[918] = 14'b000000000_0000;
storage1[919] = 14'b000000000_0000;
storage1[920] = 14'b000000101_0000;
storage1[921] = 14'b000000011_0000;
storage1[922] = 14'b000000011_0000;
storage1[923] = 14'b000000011_0000;
storage1[924] = 14'b000000011_0000;
storage1[925] = 14'b000000011_0000;
storage1[926] = 14'b000000101_0000;
storage1[927] = 14'b000000101_0000;
storage1[928] = 14'b000000011_0000;
storage1[929] = 14'b000000011_0000;
storage1[930] = 14'b000000101_0000;
storage1[931] = 14'b000000011_0000;
storage1[932] = 14'b000000101_0000;
storage1[933] = 14'b000000101_0000;
storage1[934] = 14'b000000101_0000;
storage1[935] = 14'b000000101_0000;
storage1[936] = 14'b000000101_0000;
storage1[937] = 14'b000000011_0000;
storage1[938] = 14'b000000101_0000;
storage1[939] = 14'b000000110_0000;
storage1[940] = 14'b000000101_0000;
storage1[941] = 14'b000000101_0000;
storage1[942] = 14'b000000101_0000;
storage1[943] = 14'b000000101_0000;
storage1[944] = 14'b000000101_0000;
storage1[945] = 14'b000000110_0000;
storage1[946] = 14'b000000101_0000;
storage1[947] = 14'b000000101_0000;
storage1[948] = 14'b000000101_0000;
storage1[949] = 14'b000000010_0000;
storage1[950] = 14'b000000001_0000;
storage1[951] = 14'b000000001_0000;
storage1[952] = 14'b000000000_0000;
storage1[953] = 14'b000000000_0000;
storage1[954] = 14'b000000001_0000;
storage1[955] = 14'b000000001_0000;
storage1[956] = 14'b000000001_0000;
storage1[957] = 14'b000000001_0000;
storage1[958] = 14'b000000000_0000;
storage1[959] = 14'b000000001_0000;
storage1[960] = 14'b000000101_0000;
storage1[961] = 14'b000000011_0000;
storage1[962] = 14'b000000010_0000;
storage1[963] = 14'b000000010_0000;
storage1[964] = 14'b000000010_0000;
storage1[965] = 14'b000000010_0000;
storage1[966] = 14'b000000011_0000;
storage1[967] = 14'b000000101_0000;
storage1[968] = 14'b000000101_0000;
storage1[969] = 14'b000000010_0000;
storage1[970] = 14'b000000010_0000;
storage1[971] = 14'b000000011_0000;
storage1[972] = 14'b000000011_0000;
storage1[973] = 14'b000000101_0000;
storage1[974] = 14'b000000101_0000;
storage1[975] = 14'b000000110_0000;
storage1[976] = 14'b000001001_0000;
storage1[977] = 14'b000000111_0000;
storage1[978] = 14'b000000101_0000;
storage1[979] = 14'b000000110_0000;
storage1[980] = 14'b000000101_0000;
storage1[981] = 14'b000000101_0000;
storage1[982] = 14'b000000010_0000;
storage1[983] = 14'b000000010_0000;
storage1[984] = 14'b000000010_0000;
storage1[985] = 14'b000000011_0000;
storage1[986] = 14'b000000101_0000;
storage1[987] = 14'b000000101_0000;
storage1[988] = 14'b000000110_0000;
storage1[989] = 14'b000000010_0000;
storage1[990] = 14'b000000001_0000;
storage1[991] = 14'b000000001_0000;
storage1[992] = 14'b000000001_0000;
storage1[993] = 14'b000000001_0000;
storage1[994] = 14'b000000001_0000;
storage1[995] = 14'b000000001_0000;
storage1[996] = 14'b000000001_0000;
storage1[997] = 14'b000000000_0000;
storage1[998] = 14'b000000001_0000;
storage1[999] = 14'b000000000_0000;
storage1[1000] = 14'b000000101_0000;
storage1[1001] = 14'b000000101_0000;
storage1[1002] = 14'b000000011_0000;
storage1[1003] = 14'b000000001_0000;
storage1[1004] = 14'b000000000_0000;
storage1[1005] = 14'b000000001_0000;
storage1[1006] = 14'b000000011_0000;
storage1[1007] = 14'b000000011_0000;
storage1[1008] = 14'b000000010_0000;
storage1[1009] = 14'b000000001_0000;
storage1[1010] = 14'b000000010_0000;
storage1[1011] = 14'b000000010_0000;
storage1[1012] = 14'b000000101_0000;
storage1[1013] = 14'b000000101_0000;
storage1[1014] = 14'b000000101_0000;
storage1[1015] = 14'b000000111_0000;
storage1[1016] = 14'b000011000_0000;
storage1[1017] = 14'b000110110_0000;
storage1[1018] = 14'b000000011_0000;
storage1[1019] = 14'b000000101_0000;
storage1[1020] = 14'b000000011_0000;
storage1[1021] = 14'b000000011_0000;
storage1[1022] = 14'b000000001_0000;
storage1[1023] = 14'b000000001_0000;
storage1[1024] = 14'b000000001_0000;
storage1[1025] = 14'b000000010_0000;
storage1[1026] = 14'b000000101_0000;
storage1[1027] = 14'b000000101_0000;
storage1[1028] = 14'b000000110_0000;
storage1[1029] = 14'b000000010_0000;
storage1[1030] = 14'b000000001_0000;
storage1[1031] = 14'b000000001_0000;
storage1[1032] = 14'b000000001_0000;
storage1[1033] = 14'b000000001_0000;
storage1[1034] = 14'b000000000_0000;
storage1[1035] = 14'b000000001_0000;
storage1[1036] = 14'b000000001_0000;
storage1[1037] = 14'b000000001_0000;
storage1[1038] = 14'b000000000_0000;
storage1[1039] = 14'b000000001_0000;
storage1[1040] = 14'b000000011_0000;
storage1[1041] = 14'b000000011_0000;
storage1[1042] = 14'b000000101_0000;
storage1[1043] = 14'b000000010_0000;
storage1[1044] = 14'b000000001_0000;
storage1[1045] = 14'b000000001_0000;
storage1[1046] = 14'b000000101_0000;
storage1[1047] = 14'b000000101_0000;
storage1[1048] = 14'b000000010_0000;
storage1[1049] = 14'b000000001_0000;
storage1[1050] = 14'b000000010_0000;
storage1[1051] = 14'b000000011_0000;
storage1[1052] = 14'b000000101_0000;
storage1[1053] = 14'b000000101_0000;
storage1[1054] = 14'b000000101_0000;
storage1[1055] = 14'b000000101_0000;
storage1[1056] = 14'b000010000_0000;
storage1[1057] = 14'b000111101_0000;
storage1[1058] = 14'b000000101_0000;
storage1[1059] = 14'b000000101_0000;
storage1[1060] = 14'b000000101_0000;
storage1[1061] = 14'b000000011_0000;
storage1[1062] = 14'b000000001_0000;
storage1[1063] = 14'b000000010_0000;
storage1[1064] = 14'b000000001_0000;
storage1[1065] = 14'b000000010_0000;
storage1[1066] = 14'b000000110_0000;
storage1[1067] = 14'b000000101_0000;
storage1[1068] = 14'b000000101_0000;
storage1[1069] = 14'b000000010_0000;
storage1[1070] = 14'b000000001_0000;
storage1[1071] = 14'b000000001_0000;
storage1[1072] = 14'b000000001_0000;
storage1[1073] = 14'b000000010_0000;
storage1[1074] = 14'b000000001_0000;
storage1[1075] = 14'b000000010_0000;
storage1[1076] = 14'b000000001_0000;
storage1[1077] = 14'b000000000_0000;
storage1[1078] = 14'b000000000_0000;
storage1[1079] = 14'b000000001_0000;
storage1[1080] = 14'b000000101_0000;
storage1[1081] = 14'b000000101_0000;
storage1[1082] = 14'b000000011_0000;
storage1[1083] = 14'b000000011_0000;
storage1[1084] = 14'b000000011_0000;
storage1[1085] = 14'b000000010_0000;
storage1[1086] = 14'b000000011_0000;
storage1[1087] = 14'b000000011_0000;
storage1[1088] = 14'b000000010_0000;
storage1[1089] = 14'b000000011_0000;
storage1[1090] = 14'b000000101_0000;
storage1[1091] = 14'b000000101_0000;
storage1[1092] = 14'b000000101_0000;
storage1[1093] = 14'b000000101_0000;
storage1[1094] = 14'b000000011_0000;
storage1[1095] = 14'b000000110_0000;
storage1[1096] = 14'b000000101_0000;
storage1[1097] = 14'b000000101_0000;
storage1[1098] = 14'b000000101_0000;
storage1[1099] = 14'b000000101_0000;
storage1[1100] = 14'b000000101_0000;
storage1[1101] = 14'b000000101_0000;
storage1[1102] = 14'b000000101_0000;
storage1[1103] = 14'b000000101_0000;
storage1[1104] = 14'b000000101_0000;
storage1[1105] = 14'b000000101_0000;
storage1[1106] = 14'b000000101_0000;
storage1[1107] = 14'b000000101_0000;
storage1[1108] = 14'b000000101_0000;
storage1[1109] = 14'b000000001_0000;
storage1[1110] = 14'b000000001_0000;
storage1[1111] = 14'b000000001_0000;
storage1[1112] = 14'b000000101_0000;
storage1[1113] = 14'b000000001_0000;
storage1[1114] = 14'b000000001_0000;
storage1[1115] = 14'b000000001_0000;
storage1[1116] = 14'b000000000_0000;
storage1[1117] = 14'b000000000_0000;
storage1[1118] = 14'b000000001_0000;
storage1[1119] = 14'b000000001_0000;
storage1[1120] = 14'b000000011_0000;
storage1[1121] = 14'b000000101_0000;
storage1[1122] = 14'b000000101_0000;
storage1[1123] = 14'b000000101_0000;
storage1[1124] = 14'b000000011_0000;
storage1[1125] = 14'b000000011_0000;
storage1[1126] = 14'b000000101_0000;
storage1[1127] = 14'b000000101_0000;
storage1[1128] = 14'b000000011_0000;
storage1[1129] = 14'b000000101_0000;
storage1[1130] = 14'b000000101_0000;
storage1[1131] = 14'b000000101_0000;
storage1[1132] = 14'b000000101_0000;
storage1[1133] = 14'b000000101_0000;
storage1[1134] = 14'b000000011_0000;
storage1[1135] = 14'b000000011_0000;
storage1[1136] = 14'b000000101_0000;
storage1[1137] = 14'b000000101_0000;
storage1[1138] = 14'b000000101_0000;
storage1[1139] = 14'b000000101_0000;
storage1[1140] = 14'b000000101_0000;
storage1[1141] = 14'b000000101_0000;
storage1[1142] = 14'b000000101_0000;
storage1[1143] = 14'b000000101_0000;
storage1[1144] = 14'b000000101_0000;
storage1[1145] = 14'b000000101_0000;
storage1[1146] = 14'b000000101_0000;
storage1[1147] = 14'b000000101_0000;
storage1[1148] = 14'b000000101_0000;
storage1[1149] = 14'b000000010_0000;
storage1[1150] = 14'b000000001_0000;
storage1[1151] = 14'b000000001_0000;
storage1[1152] = 14'b000000011_0000;
storage1[1153] = 14'b000000001_0000;
storage1[1154] = 14'b000000001_0000;
storage1[1155] = 14'b000000001_0000;
storage1[1156] = 14'b000000001_0000;
storage1[1157] = 14'b000000000_0000;
storage1[1158] = 14'b000000001_0000;
storage1[1159] = 14'b000000001_0000;
storage1[1160] = 14'b000000011_0000;
storage1[1161] = 14'b000000011_0000;
storage1[1162] = 14'b000000011_0000;
storage1[1163] = 14'b000000001_0000;
storage1[1164] = 14'b000000000_0000;
storage1[1165] = 14'b000000001_0000;
storage1[1166] = 14'b000000101_0000;
storage1[1167] = 14'b000000101_0000;
storage1[1168] = 14'b000000010_0000;
storage1[1169] = 14'b000000001_0000;
storage1[1170] = 14'b000000001_0000;
storage1[1171] = 14'b000000011_0000;
storage1[1172] = 14'b000000101_0000;
storage1[1173] = 14'b000000101_0000;
storage1[1174] = 14'b000000011_0000;
storage1[1175] = 14'b000000001_0000;
storage1[1176] = 14'b000000000_0000;
storage1[1177] = 14'b000000001_0000;
storage1[1178] = 14'b000000011_0000;
storage1[1179] = 14'b000000110_0000;
storage1[1180] = 14'b000000101_0000;
storage1[1181] = 14'b000000011_0000;
storage1[1182] = 14'b000000001_0000;
storage1[1183] = 14'b000000000_0000;
storage1[1184] = 14'b000000001_0000;
storage1[1185] = 14'b000000010_0000;
storage1[1186] = 14'b000000101_0000;
storage1[1187] = 14'b000000110_0000;
storage1[1188] = 14'b000000101_0000;
storage1[1189] = 14'b000000001_0000;
storage1[1190] = 14'b000000001_0000;
storage1[1191] = 14'b000000001_0000;
storage1[1192] = 14'b000000001_0000;
storage1[1193] = 14'b000000001_0000;
storage1[1194] = 14'b000000001_0000;
storage1[1195] = 14'b000000001_0000;
storage1[1196] = 14'b000000001_0000;
storage1[1197] = 14'b000000001_0000;
storage1[1198] = 14'b000000000_0000;
storage1[1199] = 14'b000000000_0000;
storage1[1200] = 14'b000000101_0000;
storage1[1201] = 14'b000000010_0000;
storage1[1202] = 14'b000000010_0000;
storage1[1203] = 14'b000000000_0000;
storage1[1204] = 14'b000000001_0000;
storage1[1205] = 14'b000000001_0000;
storage1[1206] = 14'b000000101_0000;
storage1[1207] = 14'b000000011_0000;
storage1[1208] = 14'b000000010_0000;
storage1[1209] = 14'b000000001_0000;
storage1[1210] = 14'b000000000_0000;
storage1[1211] = 14'b000000010_0000;
storage1[1212] = 14'b000000101_0000;
storage1[1213] = 14'b000000101_0000;
storage1[1214] = 14'b000000010_0000;
storage1[1215] = 14'b000000001_0000;
storage1[1216] = 14'b000000001_0000;
storage1[1217] = 14'b000000001_0000;
storage1[1218] = 14'b000000011_0000;
storage1[1219] = 14'b000000101_0000;
storage1[1220] = 14'b000000101_0000;
storage1[1221] = 14'b000000011_0000;
storage1[1222] = 14'b000000001_0000;
storage1[1223] = 14'b000000001_0000;
storage1[1224] = 14'b000000000_0000;
storage1[1225] = 14'b000000010_0000;
storage1[1226] = 14'b000000101_0000;
storage1[1227] = 14'b000000101_0000;
storage1[1228] = 14'b000000101_0000;
storage1[1229] = 14'b000000001_0000;
storage1[1230] = 14'b000000001_0000;
storage1[1231] = 14'b000000001_0000;
storage1[1232] = 14'b000000010_0000;
storage1[1233] = 14'b000000001_0000;
storage1[1234] = 14'b000000001_0000;
storage1[1235] = 14'b000000000_0000;
storage1[1236] = 14'b000000001_0000;
storage1[1237] = 14'b000000001_0000;
storage1[1238] = 14'b000000000_0000;
storage1[1239] = 14'b000000000_0000;
storage1[1240] = 14'b000000011_0000;
storage1[1241] = 14'b000000011_0000;
storage1[1242] = 14'b000000011_0000;
storage1[1243] = 14'b000000010_0000;
storage1[1244] = 14'b000000011_0000;
storage1[1245] = 14'b000000010_0000;
storage1[1246] = 14'b000000101_0000;
storage1[1247] = 14'b000000101_0000;
storage1[1248] = 14'b000000101_0000;
storage1[1249] = 14'b000000101_0000;
storage1[1250] = 14'b000000010_0000;
storage1[1251] = 14'b000000010_0000;
storage1[1252] = 14'b000000101_0000;
storage1[1253] = 14'b000000101_0000;
storage1[1254] = 14'b000000010_0000;
storage1[1255] = 14'b000000101_0000;
storage1[1256] = 14'b000000101_0000;
storage1[1257] = 14'b000000101_0000;
storage1[1258] = 14'b000000101_0000;
storage1[1259] = 14'b000000101_0000;
storage1[1260] = 14'b000000101_0000;
storage1[1261] = 14'b000000101_0000;
storage1[1262] = 14'b000000101_0000;
storage1[1263] = 14'b000000101_0000;
storage1[1264] = 14'b000000101_0000;
storage1[1265] = 14'b000000101_0000;
storage1[1266] = 14'b000000110_0000;
storage1[1267] = 14'b000000110_0000;
storage1[1268] = 14'b000000101_0000;
storage1[1269] = 14'b000000001_0000;
storage1[1270] = 14'b000000001_0000;
storage1[1271] = 14'b000000001_0000;
storage1[1272] = 14'b000000001_0000;
storage1[1273] = 14'b000000001_0000;
storage1[1274] = 14'b000000001_0000;
storage1[1275] = 14'b000000001_0000;
storage1[1276] = 14'b000000001_0000;
storage1[1277] = 14'b000000001_0000;
storage1[1278] = 14'b000000001_0000;
storage1[1279] = 14'b000000000_0000;
storage1[1280] = 14'b000000101_0000;
storage1[1281] = 14'b000000011_0000;
storage1[1282] = 14'b000000011_0000;
storage1[1283] = 14'b000000011_0000;
storage1[1284] = 14'b000000010_0000;
storage1[1285] = 14'b000000011_0000;
storage1[1286] = 14'b000000011_0000;
storage1[1287] = 14'b000000011_0000;
storage1[1288] = 14'b000000101_0000;
storage1[1289] = 14'b000000011_0000;
storage1[1290] = 14'b000000110_0000;
storage1[1291] = 14'b000000101_0000;
storage1[1292] = 14'b000000101_0000;
storage1[1293] = 14'b000000101_0000;
storage1[1294] = 14'b000000110_0000;
storage1[1295] = 14'b000000101_0000;
storage1[1296] = 14'b000000101_0000;
storage1[1297] = 14'b000000101_0000;
storage1[1298] = 14'b000000101_0000;
storage1[1299] = 14'b000000101_0000;
storage1[1300] = 14'b000000101_0000;
storage1[1301] = 14'b000000110_0000;
storage1[1302] = 14'b000000110_0000;
storage1[1303] = 14'b000000101_0000;
storage1[1304] = 14'b000000101_0000;
storage1[1305] = 14'b000000011_0000;
storage1[1306] = 14'b000000101_0000;
storage1[1307] = 14'b000000110_0000;
storage1[1308] = 14'b000000101_0000;
storage1[1309] = 14'b000000001_0000;
storage1[1310] = 14'b000000001_0000;
storage1[1311] = 14'b000000001_0000;
storage1[1312] = 14'b000000010_0000;
storage1[1313] = 14'b000000001_0000;
storage1[1314] = 14'b000000001_0000;
storage1[1315] = 14'b000000001_0000;
storage1[1316] = 14'b000000001_0000;
storage1[1317] = 14'b000000001_0000;
storage1[1318] = 14'b000000000_0000;
storage1[1319] = 14'b000000000_0000;
storage1[1320] = 14'b000000101_0000;
storage1[1321] = 14'b000000101_0000;
storage1[1322] = 14'b000000011_0000;
storage1[1323] = 14'b000000010_0000;
storage1[1324] = 14'b000000010_0000;
storage1[1325] = 14'b000000010_0000;
storage1[1326] = 14'b000000011_0000;
storage1[1327] = 14'b000000011_0000;
storage1[1328] = 14'b000000010_0000;
storage1[1329] = 14'b000000010_0000;
storage1[1330] = 14'b000000010_0000;
storage1[1331] = 14'b000000101_0000;
storage1[1332] = 14'b000000101_0000;
storage1[1333] = 14'b000000101_0000;
storage1[1334] = 14'b000000111_0000;
storage1[1335] = 14'b000001000_0000;
storage1[1336] = 14'b000010100_0000;
storage1[1337] = 14'b000100100_0000;
storage1[1338] = 14'b000000101_0000;
storage1[1339] = 14'b000000110_0000;
storage1[1340] = 14'b000000101_0000;
storage1[1341] = 14'b000000101_0000;
storage1[1342] = 14'b000000010_0000;
storage1[1343] = 14'b000000010_0000;
storage1[1344] = 14'b000000010_0000;
storage1[1345] = 14'b000000101_0000;
storage1[1346] = 14'b000000101_0000;
storage1[1347] = 14'b000000101_0000;
storage1[1348] = 14'b000000101_0000;
storage1[1349] = 14'b000000001_0000;
storage1[1350] = 14'b000000010_0000;
storage1[1351] = 14'b000000010_0000;
storage1[1352] = 14'b000000001_0000;
storage1[1353] = 14'b000000001_0000;
storage1[1354] = 14'b000000001_0000;
storage1[1355] = 14'b000000001_0000;
storage1[1356] = 14'b000000001_0000;
storage1[1357] = 14'b000000001_0000;
storage1[1358] = 14'b000000000_0000;
storage1[1359] = 14'b000000000_0000;
storage1[1360] = 14'b000000011_0000;
storage1[1361] = 14'b000000011_0000;
storage1[1362] = 14'b000000010_0000;
storage1[1363] = 14'b000000011_0000;
storage1[1364] = 14'b000000101_0000;
storage1[1365] = 14'b000000101_0000;
storage1[1366] = 14'b000000101_0000;
storage1[1367] = 14'b000000101_0000;
storage1[1368] = 14'b000000001_0000;
storage1[1369] = 14'b000000001_0000;
storage1[1370] = 14'b000000001_0000;
storage1[1371] = 14'b000000101_0000;
storage1[1372] = 14'b000000101_0000;
storage1[1373] = 14'b000000101_0000;
storage1[1374] = 14'b000001010_0000;
storage1[1375] = 14'b000010000_0000;
storage1[1376] = 14'b000110000_0000;
storage1[1377] = 14'b001101101_0000;
storage1[1378] = 14'b000001100_0000;
storage1[1379] = 14'b000000110_0000;
storage1[1380] = 14'b000000101_0000;
storage1[1381] = 14'b000000010_0000;
storage1[1382] = 14'b000000001_0000;
storage1[1383] = 14'b000000001_0000;
storage1[1384] = 14'b000000001_0000;
storage1[1385] = 14'b000000011_0000;
storage1[1386] = 14'b000000101_0000;
storage1[1387] = 14'b000000101_0000;
storage1[1388] = 14'b000000101_0000;
storage1[1389] = 14'b000000001_0000;
storage1[1390] = 14'b000000010_0000;
storage1[1391] = 14'b000000010_0000;
storage1[1392] = 14'b000000001_0000;
storage1[1393] = 14'b000000001_0000;
storage1[1394] = 14'b000000001_0000;
storage1[1395] = 14'b000000001_0000;
storage1[1396] = 14'b000000001_0000;
storage1[1397] = 14'b000000001_0000;
storage1[1398] = 14'b000000000_0000;
storage1[1399] = 14'b000000000_0000;
storage1[1400] = 14'b000000101_0000;
storage1[1401] = 14'b000000011_0000;
storage1[1402] = 14'b000000010_0000;
storage1[1403] = 14'b000000101_0000;
storage1[1404] = 14'b000001110_0000;
storage1[1405] = 14'b000001001_0000;
storage1[1406] = 14'b000000101_0000;
storage1[1407] = 14'b000000101_0000;
storage1[1408] = 14'b000000010_0000;
storage1[1409] = 14'b000000010_0000;
storage1[1410] = 14'b000000001_0000;
storage1[1411] = 14'b000000101_0000;
storage1[1412] = 14'b000000110_0000;
storage1[1413] = 14'b000000110_0000;
storage1[1414] = 14'b000000111_0000;
storage1[1415] = 14'b000001000_0000;
storage1[1416] = 14'b000101010_0000;
storage1[1417] = 14'b001000101_0000;
storage1[1418] = 14'b000001000_0000;
storage1[1419] = 14'b000000101_0000;
storage1[1420] = 14'b000000101_0000;
storage1[1421] = 14'b000000011_0000;
storage1[1422] = 14'b000000010_0000;
storage1[1423] = 14'b000000010_0000;
storage1[1424] = 14'b000000010_0000;
storage1[1425] = 14'b000000011_0000;
storage1[1426] = 14'b000000101_0000;
storage1[1427] = 14'b000000101_0000;
storage1[1428] = 14'b000000101_0000;
storage1[1429] = 14'b000000001_0000;
storage1[1430] = 14'b000000001_0000;
storage1[1431] = 14'b000000001_0000;
storage1[1432] = 14'b000000001_0000;
storage1[1433] = 14'b000000001_0000;
storage1[1434] = 14'b000000010_0000;
storage1[1435] = 14'b000000001_0000;
storage1[1436] = 14'b000000000_0000;
storage1[1437] = 14'b000000000_0000;
storage1[1438] = 14'b000000000_0000;
storage1[1439] = 14'b000000001_0000;
storage1[1440] = 14'b000000101_0000;
storage1[1441] = 14'b000000101_0000;
storage1[1442] = 14'b000000011_0000;
storage1[1443] = 14'b000000011_0000;
storage1[1444] = 14'b000000101_0000;
storage1[1445] = 14'b000000101_0000;
storage1[1446] = 14'b000000101_0000;
storage1[1447] = 14'b000000101_0000;
storage1[1448] = 14'b000000101_0000;
storage1[1449] = 14'b000000101_0000;
storage1[1450] = 14'b000000011_0000;
storage1[1451] = 14'b000000101_0000;
storage1[1452] = 14'b000000101_0000;
storage1[1453] = 14'b000000110_0000;
storage1[1454] = 14'b000000101_0000;
storage1[1455] = 14'b000000101_0000;
storage1[1456] = 14'b000000101_0000;
storage1[1457] = 14'b000000101_0000;
storage1[1458] = 14'b000000101_0000;
storage1[1459] = 14'b000000101_0000;
storage1[1460] = 14'b000000101_0000;
storage1[1461] = 14'b000000101_0000;
storage1[1462] = 14'b000000110_0000;
storage1[1463] = 14'b000000101_0000;
storage1[1464] = 14'b000000110_0000;
storage1[1465] = 14'b000000101_0000;
storage1[1466] = 14'b000000101_0000;
storage1[1467] = 14'b000000101_0000;
storage1[1468] = 14'b000000101_0000;
storage1[1469] = 14'b000000001_0000;
storage1[1470] = 14'b000000001_0000;
storage1[1471] = 14'b000000001_0000;
storage1[1472] = 14'b000000001_0000;
storage1[1473] = 14'b000000001_0000;
storage1[1474] = 14'b000000001_0000;
storage1[1475] = 14'b000000001_0000;
storage1[1476] = 14'b000000001_0000;
storage1[1477] = 14'b000000000_0000;
storage1[1478] = 14'b000000001_0000;
storage1[1479] = 14'b000000001_0000;
storage1[1480] = 14'b000000011_0000;
storage1[1481] = 14'b000000010_0000;
storage1[1482] = 14'b000000011_0000;
storage1[1483] = 14'b000000101_0000;
storage1[1484] = 14'b000000101_0000;
storage1[1485] = 14'b000000011_0000;
storage1[1486] = 14'b000000101_0000;
storage1[1487] = 14'b000000011_0000;
storage1[1488] = 14'b000000011_0000;
storage1[1489] = 14'b000000101_0000;
storage1[1490] = 14'b000000011_0000;
storage1[1491] = 14'b000000101_0000;
storage1[1492] = 14'b000000101_0000;
storage1[1493] = 14'b000000110_0000;
storage1[1494] = 14'b000000011_0000;
storage1[1495] = 14'b000000101_0000;
storage1[1496] = 14'b000000101_0000;
storage1[1497] = 14'b000000101_0000;
storage1[1498] = 14'b000000101_0000;
storage1[1499] = 14'b000000101_0000;
storage1[1500] = 14'b000000101_0000;
storage1[1501] = 14'b000000110_0000;
storage1[1502] = 14'b000000101_0000;
storage1[1503] = 14'b000000101_0000;
storage1[1504] = 14'b000000101_0000;
storage1[1505] = 14'b000000101_0000;
storage1[1506] = 14'b000000101_0000;
storage1[1507] = 14'b000000101_0000;
storage1[1508] = 14'b000000101_0000;
storage1[1509] = 14'b000000010_0000;
storage1[1510] = 14'b000000010_0000;
storage1[1511] = 14'b000000001_0000;
storage1[1512] = 14'b000000001_0000;
storage1[1513] = 14'b000000001_0000;
storage1[1514] = 14'b000000001_0000;
storage1[1515] = 14'b000000001_0000;
storage1[1516] = 14'b000000001_0000;
storage1[1517] = 14'b000000001_0000;
storage1[1518] = 14'b000000010_0000;
storage1[1519] = 14'b000000001_0000;
storage1[1520] = 14'b000000011_0000;
storage1[1521] = 14'b000000101_0000;
storage1[1522] = 14'b000000010_0000;
storage1[1523] = 14'b000000001_0000;
storage1[1524] = 14'b000000001_0000;
storage1[1525] = 14'b000000010_0000;
storage1[1526] = 14'b000000101_0000;
storage1[1527] = 14'b000000101_0000;
storage1[1528] = 14'b000000001_0000;
storage1[1529] = 14'b000000001_0000;
storage1[1530] = 14'b000000001_0000;
storage1[1531] = 14'b000000101_0000;
storage1[1532] = 14'b000000110_0000;
storage1[1533] = 14'b000000101_0000;
storage1[1534] = 14'b000000001_0000;
storage1[1535] = 14'b000000010_0000;
storage1[1536] = 14'b000000001_0000;
storage1[1537] = 14'b000000001_0000;
storage1[1538] = 14'b000000101_0000;
storage1[1539] = 14'b000000101_0000;
storage1[1540] = 14'b000000101_0000;
storage1[1541] = 14'b000000010_0000;
storage1[1542] = 14'b000000001_0000;
storage1[1543] = 14'b000000010_0000;
storage1[1544] = 14'b000000001_0000;
storage1[1545] = 14'b000000011_0000;
storage1[1546] = 14'b000000101_0000;
storage1[1547] = 14'b000000101_0000;
storage1[1548] = 14'b000000101_0000;
storage1[1549] = 14'b000000001_0000;
storage1[1550] = 14'b000000010_0000;
storage1[1551] = 14'b000000010_0000;
storage1[1552] = 14'b000000001_0000;
storage1[1553] = 14'b000000010_0000;
storage1[1554] = 14'b000000001_0000;
storage1[1555] = 14'b000000010_0000;
storage1[1556] = 14'b000000001_0000;
storage1[1557] = 14'b000000010_0000;
storage1[1558] = 14'b000000111_0000;
storage1[1559] = 14'b000000001_0000;
storage1[1560] = 14'b000000010_0000;
storage1[1561] = 14'b000000011_0000;
storage1[1562] = 14'b000000010_0000;
storage1[1563] = 14'b000000001_0000;
storage1[1564] = 14'b000000010_0000;
storage1[1565] = 14'b000000010_0000;
storage1[1566] = 14'b000000011_0000;
storage1[1567] = 14'b000000101_0000;
storage1[1568] = 14'b000000000_0000;
storage1[1569] = 14'b000000001_0000;
storage1[1570] = 14'b000000001_0000;
storage1[1571] = 14'b000000101_0000;
storage1[1572] = 14'b000000101_0000;
storage1[1573] = 14'b000000110_0000;
storage1[1574] = 14'b000000001_0000;
storage1[1575] = 14'b000000001_0000;
storage1[1576] = 14'b000000001_0000;
storage1[1577] = 14'b000000001_0000;
storage1[1578] = 14'b000000101_0000;
storage1[1579] = 14'b000000110_0000;
storage1[1580] = 14'b000000110_0000;
storage1[1581] = 14'b000000010_0000;
storage1[1582] = 14'b000000001_0000;
storage1[1583] = 14'b000000010_0000;
storage1[1584] = 14'b000000001_0000;
storage1[1585] = 14'b000000101_0000;
storage1[1586] = 14'b000000101_0000;
storage1[1587] = 14'b000000101_0000;
storage1[1588] = 14'b000000101_0000;
storage1[1589] = 14'b000000001_0000;
storage1[1590] = 14'b000000001_0000;
storage1[1591] = 14'b000000001_0000;
storage1[1592] = 14'b000000010_0000;
storage1[1593] = 14'b000000010_0000;
storage1[1594] = 14'b000000001_0000;
storage1[1595] = 14'b000000001_0000;
storage1[1596] = 14'b000000001_0000;
storage1[1597] = 14'b000000001_0000;
storage1[1598] = 14'b000000001_0000;
storage1[1599] = 14'b000000001_0000;
// image 2
storage1[1600] = 14'b001100100_0000;
storage1[1601] = 14'b001101000_0000;
storage1[1602] = 14'b001100101_0000;
storage1[1603] = 14'b001101011_0000;
storage1[1604] = 14'b001101101_0000;
storage1[1605] = 14'b001110001_0000;
storage1[1606] = 14'b001110101_0000;
storage1[1607] = 14'b001111001_0000;
storage1[1608] = 14'b001111111_0000;
storage1[1609] = 14'b010000011_0000;
storage1[1610] = 14'b010000110_0000;
storage1[1611] = 14'b010001101_0000;
storage1[1612] = 14'b010001111_0000;
storage1[1613] = 14'b010010011_0000;
storage1[1614] = 14'b010010101_0000;
storage1[1615] = 14'b010010011_0000;
storage1[1616] = 14'b010010111_0000;
storage1[1617] = 14'b010010110_0000;
storage1[1618] = 14'b010010010_0000;
storage1[1619] = 14'b010010000_0000;
storage1[1620] = 14'b010001111_0000;
storage1[1621] = 14'b010001101_0000;
storage1[1622] = 14'b010001101_0000;
storage1[1623] = 14'b010001011_0000;
storage1[1624] = 14'b010001000_0000;
storage1[1625] = 14'b010000100_0000;
storage1[1626] = 14'b010110110_0000;
storage1[1627] = 14'b011101101_0000;
storage1[1628] = 14'b010001111_0000;
storage1[1629] = 14'b010000000_0000;
storage1[1630] = 14'b010000001_0000;
storage1[1631] = 14'b001111110_0000;
storage1[1632] = 14'b001111110_0000;
storage1[1633] = 14'b010000000_0000;
storage1[1634] = 14'b001111111_0000;
storage1[1635] = 14'b001111111_0000;
storage1[1636] = 14'b001111101_0000;
storage1[1637] = 14'b001111101_0000;
storage1[1638] = 14'b001111100_0000;
storage1[1639] = 14'b001111100_0000;
storage1[1640] = 14'b001011011_0000;
storage1[1641] = 14'b001100001_0000;
storage1[1642] = 14'b001011111_0000;
storage1[1643] = 14'b001100100_0000;
storage1[1644] = 14'b001101000_0000;
storage1[1645] = 14'b001101000_0000;
storage1[1646] = 14'b001101100_0000;
storage1[1647] = 14'b001110000_0000;
storage1[1648] = 14'b001110010_0000;
storage1[1649] = 14'b001110111_0000;
storage1[1650] = 14'b001111000_0000;
storage1[1651] = 14'b001111011_0000;
storage1[1652] = 14'b001111011_0000;
storage1[1653] = 14'b001111111_0000;
storage1[1654] = 14'b010000001_0000;
storage1[1655] = 14'b010000010_0000;
storage1[1656] = 14'b010000010_0000;
storage1[1657] = 14'b010000001_0000;
storage1[1658] = 14'b010000000_0000;
storage1[1659] = 14'b001111111_0000;
storage1[1660] = 14'b001111111_0000;
storage1[1661] = 14'b001111110_0000;
storage1[1662] = 14'b001111101_0000;
storage1[1663] = 14'b001111100_0000;
storage1[1664] = 14'b001111101_0000;
storage1[1665] = 14'b001110110_0000;
storage1[1666] = 14'b001111011_0000;
storage1[1667] = 14'b010000110_0000;
storage1[1668] = 14'b001111001_0000;
storage1[1669] = 14'b001111000_0000;
storage1[1670] = 14'b001111111_0000;
storage1[1671] = 14'b001111111_0000;
storage1[1672] = 14'b001111110_0000;
storage1[1673] = 14'b001111110_0000;
storage1[1674] = 14'b001111111_0000;
storage1[1675] = 14'b001111101_0000;
storage1[1676] = 14'b001111110_0000;
storage1[1677] = 14'b001111101_0000;
storage1[1678] = 14'b001111110_0000;
storage1[1679] = 14'b001111110_0000;
storage1[1680] = 14'b010101101_0000;
storage1[1681] = 14'b010101101_0000;
storage1[1682] = 14'b010101110_0000;
storage1[1683] = 14'b010110001_0000;
storage1[1684] = 14'b010110010_0000;
storage1[1685] = 14'b010110111_0000;
storage1[1686] = 14'b010111010_0000;
storage1[1687] = 14'b010111001_0000;
storage1[1688] = 14'b010111100_0000;
storage1[1689] = 14'b010111110_0000;
storage1[1690] = 14'b010111111_0000;
storage1[1691] = 14'b011000001_0000;
storage1[1692] = 14'b011000011_0000;
storage1[1693] = 14'b011000011_0000;
storage1[1694] = 14'b011000110_0000;
storage1[1695] = 14'b011000110_0000;
storage1[1696] = 14'b011000110_0000;
storage1[1697] = 14'b011001001_0000;
storage1[1698] = 14'b011000111_0000;
storage1[1699] = 14'b011001001_0000;
storage1[1700] = 14'b011001000_0000;
storage1[1701] = 14'b011000111_0000;
storage1[1702] = 14'b011000110_0000;
storage1[1703] = 14'b011000101_0000;
storage1[1704] = 14'b011000101_0000;
storage1[1705] = 14'b011000110_0000;
storage1[1706] = 14'b011001001_0000;
storage1[1707] = 14'b011000111_0000;
storage1[1708] = 14'b011001001_0000;
storage1[1709] = 14'b011001001_0000;
storage1[1710] = 14'b010100100_0000;
storage1[1711] = 14'b001111101_0000;
storage1[1712] = 14'b001111101_0000;
storage1[1713] = 14'b010000000_0000;
storage1[1714] = 14'b001111111_0000;
storage1[1715] = 14'b001111111_0000;
storage1[1716] = 14'b001111110_0000;
storage1[1717] = 14'b001111111_0000;
storage1[1718] = 14'b001111110_0000;
storage1[1719] = 14'b001111101_0000;
storage1[1720] = 14'b010111010_0000;
storage1[1721] = 14'b010111010_0000;
storage1[1722] = 14'b010111000_0000;
storage1[1723] = 14'b010111010_0000;
storage1[1724] = 14'b010111100_0000;
storage1[1725] = 14'b010111110_0000;
storage1[1726] = 14'b010111110_0000;
storage1[1727] = 14'b010111111_0000;
storage1[1728] = 14'b010111111_0000;
storage1[1729] = 14'b011000010_0000;
storage1[1730] = 14'b011000010_0000;
storage1[1731] = 14'b011000010_0000;
storage1[1732] = 14'b011000101_0000;
storage1[1733] = 14'b011000011_0000;
storage1[1734] = 14'b011000110_0000;
storage1[1735] = 14'b011001000_0000;
storage1[1736] = 14'b011000111_0000;
storage1[1737] = 14'b011000101_0000;
storage1[1738] = 14'b011001000_0000;
storage1[1739] = 14'b011001000_0000;
storage1[1740] = 14'b011000111_0000;
storage1[1741] = 14'b011001000_0000;
storage1[1742] = 14'b011001000_0000;
storage1[1743] = 14'b011000101_0000;
storage1[1744] = 14'b011000011_0000;
storage1[1745] = 14'b011000100_0000;
storage1[1746] = 14'b011000110_0000;
storage1[1747] = 14'b011000100_0000;
storage1[1748] = 14'b011000110_0000;
storage1[1749] = 14'b011000110_0000;
storage1[1750] = 14'b010101111_0000;
storage1[1751] = 14'b010011101_0000;
storage1[1752] = 14'b001111101_0000;
storage1[1753] = 14'b001111111_0000;
storage1[1754] = 14'b001111111_0000;
storage1[1755] = 14'b010000000_0000;
storage1[1756] = 14'b010000001_0000;
storage1[1757] = 14'b001111110_0000;
storage1[1758] = 14'b001111110_0000;
storage1[1759] = 14'b001111110_0000;
storage1[1760] = 14'b010110111_0000;
storage1[1761] = 14'b010111010_0000;
storage1[1762] = 14'b010111000_0000;
storage1[1763] = 14'b010111100_0000;
storage1[1764] = 14'b010111101_0000;
storage1[1765] = 14'b010111100_0000;
storage1[1766] = 14'b010111101_0000;
storage1[1767] = 14'b010111110_0000;
storage1[1768] = 14'b010111111_0000;
storage1[1769] = 14'b011000011_0000;
storage1[1770] = 14'b011000000_0000;
storage1[1771] = 14'b011000001_0000;
storage1[1772] = 14'b011000011_0000;
storage1[1773] = 14'b011000110_0000;
storage1[1774] = 14'b011000110_0000;
storage1[1775] = 14'b011000110_0000;
storage1[1776] = 14'b011000110_0000;
storage1[1777] = 14'b011001001_0000;
storage1[1778] = 14'b011000111_0000;
storage1[1779] = 14'b011000111_0000;
storage1[1780] = 14'b011000110_0000;
storage1[1781] = 14'b011000111_0000;
storage1[1782] = 14'b011000111_0000;
storage1[1783] = 14'b011000110_0000;
storage1[1784] = 14'b011000110_0000;
storage1[1785] = 14'b011000101_0000;
storage1[1786] = 14'b011000111_0000;
storage1[1787] = 14'b011000101_0000;
storage1[1788] = 14'b011000110_0000;
storage1[1789] = 14'b011001011_0000;
storage1[1790] = 14'b010101111_0000;
storage1[1791] = 14'b010101100_0000;
storage1[1792] = 14'b010011000_0000;
storage1[1793] = 14'b001111111_0000;
storage1[1794] = 14'b010101100_0000;
storage1[1795] = 14'b001111010_0000;
storage1[1796] = 14'b001111111_0000;
storage1[1797] = 14'b010000000_0000;
storage1[1798] = 14'b001111110_0000;
storage1[1799] = 14'b010000000_0000;
storage1[1800] = 14'b010111111_0000;
storage1[1801] = 14'b010111100_0000;
storage1[1802] = 14'b010111010_0000;
storage1[1803] = 14'b010111111_0000;
storage1[1804] = 14'b010111111_0000;
storage1[1805] = 14'b010111110_0000;
storage1[1806] = 14'b011000010_0000;
storage1[1807] = 14'b011000000_0000;
storage1[1808] = 14'b011000001_0000;
storage1[1809] = 14'b011000011_0000;
storage1[1810] = 14'b011000101_0000;
storage1[1811] = 14'b011000110_0000;
storage1[1812] = 14'b011000101_0000;
storage1[1813] = 14'b011001000_0000;
storage1[1814] = 14'b011001001_0000;
storage1[1815] = 14'b011001100_0000;
storage1[1816] = 14'b011001011_0000;
storage1[1817] = 14'b011001011_0000;
storage1[1818] = 14'b011001011_0000;
storage1[1819] = 14'b011000111_0000;
storage1[1820] = 14'b011000111_0000;
storage1[1821] = 14'b011001001_0000;
storage1[1822] = 14'b011001001_0000;
storage1[1823] = 14'b011000111_0000;
storage1[1824] = 14'b011000111_0000;
storage1[1825] = 14'b011000110_0000;
storage1[1826] = 14'b011000111_0000;
storage1[1827] = 14'b011000110_0000;
storage1[1828] = 14'b011000110_0000;
storage1[1829] = 14'b011001001_0000;
storage1[1830] = 14'b010110000_0000;
storage1[1831] = 14'b010101101_0000;
storage1[1832] = 14'b010101001_0000;
storage1[1833] = 14'b010010101_0000;
storage1[1834] = 14'b010111110_0000;
storage1[1835] = 14'b001111100_0000;
storage1[1836] = 14'b010000001_0000;
storage1[1837] = 14'b010000000_0000;
storage1[1838] = 14'b010000001_0000;
storage1[1839] = 14'b010000000_0000;
storage1[1840] = 14'b010001111_0000;
storage1[1841] = 14'b011000001_0000;
storage1[1842] = 14'b010111111_0000;
storage1[1843] = 14'b011000001_0000;
storage1[1844] = 14'b010001100_0000;
storage1[1845] = 14'b010110000_0000;
storage1[1846] = 14'b010011000_0000;
storage1[1847] = 14'b011000101_0000;
storage1[1848] = 14'b011000100_0000;
storage1[1849] = 14'b010100010_0000;
storage1[1850] = 14'b010010011_0000;
storage1[1851] = 14'b010010101_0000;
storage1[1852] = 14'b010111001_0000;
storage1[1853] = 14'b011001001_0000;
storage1[1854] = 14'b011001010_0000;
storage1[1855] = 14'b010100001_0000;
storage1[1856] = 14'b010010010_0000;
storage1[1857] = 14'b010110101_0000;
storage1[1858] = 14'b010011101_0000;
storage1[1859] = 14'b010110110_0000;
storage1[1860] = 14'b011000111_0000;
storage1[1861] = 14'b011000110_0000;
storage1[1862] = 14'b010100001_0000;
storage1[1863] = 14'b010001000_0000;
storage1[1864] = 14'b010001100_0000;
storage1[1865] = 14'b010000111_0000;
storage1[1866] = 14'b010101110_0000;
storage1[1867] = 14'b011001000_0000;
storage1[1868] = 14'b011001010_0000;
storage1[1869] = 14'b011001010_0000;
storage1[1870] = 14'b010101000_0000;
storage1[1871] = 14'b010101101_0000;
storage1[1872] = 14'b010101001_0000;
storage1[1873] = 14'b010101000_0000;
storage1[1874] = 14'b011010100_0000;
storage1[1875] = 14'b001111101_0000;
storage1[1876] = 14'b010000010_0000;
storage1[1877] = 14'b010000010_0000;
storage1[1878] = 14'b010000000_0000;
storage1[1879] = 14'b010000001_0000;
storage1[1880] = 14'b010101111_0000;
storage1[1881] = 14'b011000100_0000;
storage1[1882] = 14'b011000000_0000;
storage1[1883] = 14'b011000000_0000;
storage1[1884] = 14'b011000001_0000;
storage1[1885] = 14'b011110000_0000;
storage1[1886] = 14'b010111111_0000;
storage1[1887] = 14'b011000011_0000;
storage1[1888] = 14'b011000111_0000;
storage1[1889] = 14'b010100100_0000;
storage1[1890] = 14'b011000100_0000;
storage1[1891] = 14'b011100110_0000;
storage1[1892] = 14'b010111110_0000;
storage1[1893] = 14'b011001011_0000;
storage1[1894] = 14'b011001011_0000;
storage1[1895] = 14'b010100000_0000;
storage1[1896] = 14'b010011101_0000;
storage1[1897] = 14'b011111001_0000;
storage1[1898] = 14'b010111110_0000;
storage1[1899] = 14'b010111000_0000;
storage1[1900] = 14'b011001000_0000;
storage1[1901] = 14'b011001000_0000;
storage1[1902] = 14'b010011101_0000;
storage1[1903] = 14'b010001010_0000;
storage1[1904] = 14'b010010101_0000;
storage1[1905] = 14'b010001001_0000;
storage1[1906] = 14'b010101110_0000;
storage1[1907] = 14'b011000111_0000;
storage1[1908] = 14'b011001001_0000;
storage1[1909] = 14'b011001100_0000;
storage1[1910] = 14'b010001001_0000;
storage1[1911] = 14'b010101101_0000;
storage1[1912] = 14'b010101011_0000;
storage1[1913] = 14'b010101001_0000;
storage1[1914] = 14'b010100111_0000;
storage1[1915] = 14'b010001111_0000;
storage1[1916] = 14'b010000010_0000;
storage1[1917] = 14'b010000011_0000;
storage1[1918] = 14'b010000001_0000;
storage1[1919] = 14'b010000001_0000;
storage1[1920] = 14'b010011101_0000;
storage1[1921] = 14'b011000011_0000;
storage1[1922] = 14'b011000100_0000;
storage1[1923] = 14'b011000011_0000;
storage1[1924] = 14'b011000011_0000;
storage1[1925] = 14'b011111011_0000;
storage1[1926] = 14'b011000111_0000;
storage1[1927] = 14'b011000110_0000;
storage1[1928] = 14'b011000110_0000;
storage1[1929] = 14'b010100011_0000;
storage1[1930] = 14'b011011001_0000;
storage1[1931] = 14'b011100110_0000;
storage1[1932] = 14'b011000100_0000;
storage1[1933] = 14'b011001001_0000;
storage1[1934] = 14'b011001011_0000;
storage1[1935] = 14'b010011010_0000;
storage1[1936] = 14'b010010111_0000;
storage1[1937] = 14'b011111001_0000;
storage1[1938] = 14'b010110100_0000;
storage1[1939] = 14'b010111011_0000;
storage1[1940] = 14'b011001010_0000;
storage1[1941] = 14'b011001010_0000;
storage1[1942] = 14'b010011101_0000;
storage1[1943] = 14'b010000000_0000;
storage1[1944] = 14'b010001000_0000;
storage1[1945] = 14'b001111110_0000;
storage1[1946] = 14'b010101101_0000;
storage1[1947] = 14'b011000111_0000;
storage1[1948] = 14'b011001011_0000;
storage1[1949] = 14'b011001000_0000;
storage1[1950] = 14'b010000111_0000;
storage1[1951] = 14'b010011011_0000;
storage1[1952] = 14'b010011111_0000;
storage1[1953] = 14'b010101001_0000;
storage1[1954] = 14'b010101001_0000;
storage1[1955] = 14'b010100101_0000;
storage1[1956] = 14'b010001100_0000;
storage1[1957] = 14'b010000011_0000;
storage1[1958] = 14'b010000100_0000;
storage1[1959] = 14'b010000011_0000;
storage1[1960] = 14'b001111010_0000;
storage1[1961] = 14'b011000011_0000;
storage1[1962] = 14'b011000101_0000;
storage1[1963] = 14'b011000100_0000;
storage1[1964] = 14'b001110001_0000;
storage1[1965] = 14'b001111110_0000;
storage1[1966] = 14'b010001011_0000;
storage1[1967] = 14'b011001011_0000;
storage1[1968] = 14'b011001011_0000;
storage1[1969] = 14'b010011000_0000;
storage1[1970] = 14'b001111010_0000;
storage1[1971] = 14'b001110100_0000;
storage1[1972] = 14'b011001100_0000;
storage1[1973] = 14'b011001100_0000;
storage1[1974] = 14'b011001101_0000;
storage1[1975] = 14'b010010110_0000;
storage1[1976] = 14'b001111111_0000;
storage1[1977] = 14'b001111101_0000;
storage1[1978] = 14'b001111010_0000;
storage1[1979] = 14'b011000011_0000;
storage1[1980] = 14'b011001101_0000;
storage1[1981] = 14'b011001011_0000;
storage1[1982] = 14'b010011111_0000;
storage1[1983] = 14'b010000001_0000;
storage1[1984] = 14'b010000000_0000;
storage1[1985] = 14'b001111110_0000;
storage1[1986] = 14'b010110011_0000;
storage1[1987] = 14'b011001110_0000;
storage1[1988] = 14'b011001100_0000;
storage1[1989] = 14'b011000101_0000;
storage1[1990] = 14'b010001001_0000;
storage1[1991] = 14'b010011001_0000;
storage1[1992] = 14'b010011111_0000;
storage1[1993] = 14'b010011101_0000;
storage1[1994] = 14'b010101011_0000;
storage1[1995] = 14'b010100101_0000;
storage1[1996] = 14'b010100001_0000;
storage1[1997] = 14'b010001100_0000;
storage1[1998] = 14'b010000100_0000;
storage1[1999] = 14'b010000011_0000;
storage1[2000] = 14'b001111100_0000;
storage1[2001] = 14'b011000010_0000;
storage1[2002] = 14'b011000101_0000;
storage1[2003] = 14'b011000010_0000;
storage1[2004] = 14'b001110001_0000;
storage1[2005] = 14'b001110110_0000;
storage1[2006] = 14'b010010001_0000;
storage1[2007] = 14'b011001000_0000;
storage1[2008] = 14'b011001000_0000;
storage1[2009] = 14'b010010010_0000;
storage1[2010] = 14'b001111001_0000;
storage1[2011] = 14'b001111000_0000;
storage1[2012] = 14'b011001111_0000;
storage1[2013] = 14'b011001100_0000;
storage1[2014] = 14'b011001110_0000;
storage1[2015] = 14'b010010000_0000;
storage1[2016] = 14'b001111111_0000;
storage1[2017] = 14'b001111110_0000;
storage1[2018] = 14'b001111101_0000;
storage1[2019] = 14'b011000101_0000;
storage1[2020] = 14'b011001101_0000;
storage1[2021] = 14'b011001001_0000;
storage1[2022] = 14'b010011011_0000;
storage1[2023] = 14'b010000011_0000;
storage1[2024] = 14'b010000100_0000;
storage1[2025] = 14'b001111110_0000;
storage1[2026] = 14'b010111001_0000;
storage1[2027] = 14'b011001011_0000;
storage1[2028] = 14'b011001011_0000;
storage1[2029] = 14'b011000110_0000;
storage1[2030] = 14'b010001101_0000;
storage1[2031] = 14'b010010111_0000;
storage1[2032] = 14'b010100111_0000;
storage1[2033] = 14'b010100000_0000;
storage1[2034] = 14'b010010010_0000;
storage1[2035] = 14'b010100110_0000;
storage1[2036] = 14'b010100110_0000;
storage1[2037] = 14'b010011110_0000;
storage1[2038] = 14'b010000011_0000;
storage1[2039] = 14'b010000100_0000;
storage1[2040] = 14'b010011010_0000;
storage1[2041] = 14'b011000000_0000;
storage1[2042] = 14'b011000011_0000;
storage1[2043] = 14'b010111100_0000;
storage1[2044] = 14'b010101111_0000;
storage1[2045] = 14'b011010100_0000;
storage1[2046] = 14'b011001101_0000;
storage1[2047] = 14'b011000111_0000;
storage1[2048] = 14'b011001001_0000;
storage1[2049] = 14'b010010100_0000;
storage1[2050] = 14'b010101111_0000;
storage1[2051] = 14'b010101010_0000;
storage1[2052] = 14'b011001111_0000;
storage1[2053] = 14'b011001111_0000;
storage1[2054] = 14'b011001110_0000;
storage1[2055] = 14'b011001000_0000;
storage1[2056] = 14'b011011011_0000;
storage1[2057] = 14'b011100011_0000;
storage1[2058] = 14'b011101001_0000;
storage1[2059] = 14'b011001011_0000;
storage1[2060] = 14'b011001101_0000;
storage1[2061] = 14'b011001110_0000;
storage1[2062] = 14'b010101011_0000;
storage1[2063] = 14'b011001011_0000;
storage1[2064] = 14'b011101000_0000;
storage1[2065] = 14'b011001111_0000;
storage1[2066] = 14'b011000011_0000;
storage1[2067] = 14'b011001110_0000;
storage1[2068] = 14'b011001110_0000;
storage1[2069] = 14'b011000100_0000;
storage1[2070] = 14'b010001011_0000;
storage1[2071] = 14'b010011000_0000;
storage1[2072] = 14'b010101000_0000;
storage1[2073] = 14'b010011110_0000;
storage1[2074] = 14'b010001110_0000;
storage1[2075] = 14'b010001110_0000;
storage1[2076] = 14'b010100101_0000;
storage1[2077] = 14'b010011101_0000;
storage1[2078] = 14'b010000011_0000;
storage1[2079] = 14'b010000101_0000;
storage1[2080] = 14'b011000101_0000;
storage1[2081] = 14'b011000011_0000;
storage1[2082] = 14'b011000100_0000;
storage1[2083] = 14'b010111001_0000;
storage1[2084] = 14'b010110110_0000;
storage1[2085] = 14'b011110011_0000;
storage1[2086] = 14'b011100010_0000;
storage1[2087] = 14'b011001000_0000;
storage1[2088] = 14'b011001001_0000;
storage1[2089] = 14'b010010110_0000;
storage1[2090] = 14'b011011110_0000;
storage1[2091] = 14'b010111110_0000;
storage1[2092] = 14'b011010000_0000;
storage1[2093] = 14'b011001101_0000;
storage1[2094] = 14'b011001110_0000;
storage1[2095] = 14'b011011111_0000;
storage1[2096] = 14'b011111001_0000;
storage1[2097] = 14'b011111001_0000;
storage1[2098] = 14'b011111010_0000;
storage1[2099] = 14'b011010000_0000;
storage1[2100] = 14'b011010000_0000;
storage1[2101] = 14'b011001111_0000;
storage1[2102] = 14'b010101010_0000;
storage1[2103] = 14'b011110010_0000;
storage1[2104] = 14'b011111100_0000;
storage1[2105] = 14'b011101100_0000;
storage1[2106] = 14'b011000011_0000;
storage1[2107] = 14'b011001100_0000;
storage1[2108] = 14'b011001101_0000;
storage1[2109] = 14'b011000011_0000;
storage1[2110] = 14'b010001001_0000;
storage1[2111] = 14'b010010100_0000;
storage1[2112] = 14'b010100001_0000;
storage1[2113] = 14'b010010100_0000;
storage1[2114] = 14'b010001111_0000;
storage1[2115] = 14'b010000101_0000;
storage1[2116] = 14'b010010101_0000;
storage1[2117] = 14'b010011111_0000;
storage1[2118] = 14'b010000101_0000;
storage1[2119] = 14'b010000110_0000;
storage1[2120] = 14'b011000011_0000;
storage1[2121] = 14'b011000110_0000;
storage1[2122] = 14'b011000101_0000;
storage1[2123] = 14'b010111110_0000;
storage1[2124] = 14'b010110011_0000;
storage1[2125] = 14'b011001001_0000;
storage1[2126] = 14'b011001010_0000;
storage1[2127] = 14'b011000111_0000;
storage1[2128] = 14'b011001001_0000;
storage1[2129] = 14'b010101010_0000;
storage1[2130] = 14'b011010011_0000;
storage1[2131] = 14'b010111101_0000;
storage1[2132] = 14'b011010001_0000;
storage1[2133] = 14'b011001101_0000;
storage1[2134] = 14'b011010001_0000;
storage1[2135] = 14'b011001111_0000;
storage1[2136] = 14'b011011110_0000;
storage1[2137] = 14'b011011000_0000;
storage1[2138] = 14'b011100001_0000;
storage1[2139] = 14'b011001011_0000;
storage1[2140] = 14'b011001101_0000;
storage1[2141] = 14'b011010000_0000;
storage1[2142] = 14'b010110011_0000;
storage1[2143] = 14'b011010001_0000;
storage1[2144] = 14'b011011011_0000;
storage1[2145] = 14'b011010101_0000;
storage1[2146] = 14'b011001010_0000;
storage1[2147] = 14'b011010000_0000;
storage1[2148] = 14'b011010000_0000;
storage1[2149] = 14'b011000101_0000;
storage1[2150] = 14'b010001001_0000;
storage1[2151] = 14'b010001100_0000;
storage1[2152] = 14'b010011111_0000;
storage1[2153] = 14'b010010001_0000;
storage1[2154] = 14'b010010011_0000;
storage1[2155] = 14'b010001001_0000;
storage1[2156] = 14'b010000111_0000;
storage1[2157] = 14'b010010011_0000;
storage1[2158] = 14'b010000111_0000;
storage1[2159] = 14'b010001000_0000;
storage1[2160] = 14'b011000110_0000;
storage1[2161] = 14'b011000100_0000;
storage1[2162] = 14'b011000110_0000;
storage1[2163] = 14'b011000010_0000;
storage1[2164] = 14'b011001001_0000;
storage1[2165] = 14'b011001010_0000;
storage1[2166] = 14'b011001000_0000;
storage1[2167] = 14'b011001000_0000;
storage1[2168] = 14'b011001001_0000;
storage1[2169] = 14'b011000101_0000;
storage1[2170] = 14'b011001100_0000;
storage1[2171] = 14'b011001100_0000;
storage1[2172] = 14'b011010010_0000;
storage1[2173] = 14'b011001111_0000;
storage1[2174] = 14'b011010000_0000;
storage1[2175] = 14'b011001110_0000;
storage1[2176] = 14'b011001101_0000;
storage1[2177] = 14'b011010000_0000;
storage1[2178] = 14'b011001100_0000;
storage1[2179] = 14'b011001111_0000;
storage1[2180] = 14'b011010000_0000;
storage1[2181] = 14'b011010000_0000;
storage1[2182] = 14'b010111111_0000;
storage1[2183] = 14'b011001110_0000;
storage1[2184] = 14'b011001101_0000;
storage1[2185] = 14'b011001111_0000;
storage1[2186] = 14'b011001011_0000;
storage1[2187] = 14'b011001110_0000;
storage1[2188] = 14'b011001110_0000;
storage1[2189] = 14'b011000011_0000;
storage1[2190] = 14'b010101001_0000;
storage1[2191] = 14'b010001100_0000;
storage1[2192] = 14'b010011110_0000;
storage1[2193] = 14'b010010010_0000;
storage1[2194] = 14'b010001111_0000;
storage1[2195] = 14'b010001011_0000;
storage1[2196] = 14'b010001001_0000;
storage1[2197] = 14'b010010001_0000;
storage1[2198] = 14'b010001011_0000;
storage1[2199] = 14'b010001011_0000;
storage1[2200] = 14'b010110111_0000;
storage1[2201] = 14'b010111111_0000;
storage1[2202] = 14'b010111111_0000;
storage1[2203] = 14'b010111010_0000;
storage1[2204] = 14'b010110110_0000;
storage1[2205] = 14'b010110111_0000;
storage1[2206] = 14'b010111100_0000;
storage1[2207] = 14'b011000011_0000;
storage1[2208] = 14'b011000011_0000;
storage1[2209] = 14'b010111000_0000;
storage1[2210] = 14'b010111111_0000;
storage1[2211] = 14'b010111111_0000;
storage1[2212] = 14'b011001010_0000;
storage1[2213] = 14'b011001101_0000;
storage1[2214] = 14'b011001001_0000;
storage1[2215] = 14'b011001011_0000;
storage1[2216] = 14'b011010101_0000;
storage1[2217] = 14'b011001011_0000;
storage1[2218] = 14'b011000100_0000;
storage1[2219] = 14'b011001011_0000;
storage1[2220] = 14'b011001100_0000;
storage1[2221] = 14'b011010001_0000;
storage1[2222] = 14'b010110111_0000;
storage1[2223] = 14'b010111101_0000;
storage1[2224] = 14'b010111101_0000;
storage1[2225] = 14'b010111100_0000;
storage1[2226] = 14'b011001101_0000;
storage1[2227] = 14'b011010000_0000;
storage1[2228] = 14'b011010000_0000;
storage1[2229] = 14'b010111110_0000;
storage1[2230] = 14'b010100100_0000;
storage1[2231] = 14'b010100011_0000;
storage1[2232] = 14'b010011001_0000;
storage1[2233] = 14'b010010010_0000;
storage1[2234] = 14'b010010000_0000;
storage1[2235] = 14'b010001000_0000;
storage1[2236] = 14'b010001011_0000;
storage1[2237] = 14'b010010100_0000;
storage1[2238] = 14'b010001101_0000;
storage1[2239] = 14'b010001100_0000;
storage1[2240] = 14'b010110000_0000;
storage1[2241] = 14'b011000111_0000;
storage1[2242] = 14'b011001000_0000;
storage1[2243] = 14'b010101110_0000;
storage1[2244] = 14'b010010101_0000;
storage1[2245] = 14'b010011110_0000;
storage1[2246] = 14'b010111000_0000;
storage1[2247] = 14'b011001000_0000;
storage1[2248] = 14'b011001100_0000;
storage1[2249] = 14'b010001100_0000;
storage1[2250] = 14'b010100111_0000;
storage1[2251] = 14'b010100101_0000;
storage1[2252] = 14'b011010001_0000;
storage1[2253] = 14'b011010001_0000;
storage1[2254] = 14'b011010001_0000;
storage1[2255] = 14'b011111011_0000;
storage1[2256] = 14'b011111100_0000;
storage1[2257] = 14'b011110111_0000;
storage1[2258] = 14'b011001010_0000;
storage1[2259] = 14'b011010010_0000;
storage1[2260] = 14'b011010010_0000;
storage1[2261] = 14'b011010011_0000;
storage1[2262] = 14'b010010100_0000;
storage1[2263] = 14'b010110001_0000;
storage1[2264] = 14'b010101001_0000;
storage1[2265] = 14'b010100011_0000;
storage1[2266] = 14'b011010110_0000;
storage1[2267] = 14'b011010010_0000;
storage1[2268] = 14'b011010010_0000;
storage1[2269] = 14'b011000001_0000;
storage1[2270] = 14'b010011010_0000;
storage1[2271] = 14'b010100000_0000;
storage1[2272] = 14'b010100111_0000;
storage1[2273] = 14'b010010110_0000;
storage1[2274] = 14'b010001101_0000;
storage1[2275] = 14'b010000111_0000;
storage1[2276] = 14'b010001101_0000;
storage1[2277] = 14'b010010101_0000;
storage1[2278] = 14'b010001110_0000;
storage1[2279] = 14'b010001101_0000;
storage1[2280] = 14'b010101110_0000;
storage1[2281] = 14'b011001000_0000;
storage1[2282] = 14'b011001010_0000;
storage1[2283] = 14'b010101101_0000;
storage1[2284] = 14'b010001110_0000;
storage1[2285] = 14'b010001111_0000;
storage1[2286] = 14'b010110110_0000;
storage1[2287] = 14'b011001010_0000;
storage1[2288] = 14'b011001110_0000;
storage1[2289] = 14'b010001011_0000;
storage1[2290] = 14'b010010101_0000;
storage1[2291] = 14'b010011111_0000;
storage1[2292] = 14'b011010001_0000;
storage1[2293] = 14'b011010010_0000;
storage1[2294] = 14'b011010010_0000;
storage1[2295] = 14'b011101001_0000;
storage1[2296] = 14'b011110111_0000;
storage1[2297] = 14'b011101100_0000;
storage1[2298] = 14'b010111110_0000;
storage1[2299] = 14'b011010001_0000;
storage1[2300] = 14'b011010011_0000;
storage1[2301] = 14'b011010110_0000;
storage1[2302] = 14'b010010101_0000;
storage1[2303] = 14'b010100100_0000;
storage1[2304] = 14'b010100011_0000;
storage1[2305] = 14'b010011011_0000;
storage1[2306] = 14'b011010111_0000;
storage1[2307] = 14'b011010011_0000;
storage1[2308] = 14'b011010010_0000;
storage1[2309] = 14'b010111111_0000;
storage1[2310] = 14'b010010100_0000;
storage1[2311] = 14'b010011100_0000;
storage1[2312] = 14'b010011110_0000;
storage1[2313] = 14'b010101000_0000;
storage1[2314] = 14'b010010011_0000;
storage1[2315] = 14'b010000101_0000;
storage1[2316] = 14'b010001100_0000;
storage1[2317] = 14'b010011011_0000;
storage1[2318] = 14'b010001111_0000;
storage1[2319] = 14'b010001110_0000;
storage1[2320] = 14'b011000111_0000;
storage1[2321] = 14'b011000110_0000;
storage1[2322] = 14'b011000100_0000;
storage1[2323] = 14'b011000110_0000;
storage1[2324] = 14'b011001101_0000;
storage1[2325] = 14'b011001110_0000;
storage1[2326] = 14'b011001000_0000;
storage1[2327] = 14'b011001010_0000;
storage1[2328] = 14'b011001001_0000;
storage1[2329] = 14'b011001101_0000;
storage1[2330] = 14'b011001111_0000;
storage1[2331] = 14'b011001101_0000;
storage1[2332] = 14'b011010001_0000;
storage1[2333] = 14'b011001111_0000;
storage1[2334] = 14'b011001100_0000;
storage1[2335] = 14'b011001111_0000;
storage1[2336] = 14'b011010000_0000;
storage1[2337] = 14'b011001110_0000;
storage1[2338] = 14'b011001111_0000;
storage1[2339] = 14'b011010011_0000;
storage1[2340] = 14'b011010010_0000;
storage1[2341] = 14'b011010000_0000;
storage1[2342] = 14'b011001110_0000;
storage1[2343] = 14'b011010010_0000;
storage1[2344] = 14'b011010010_0000;
storage1[2345] = 14'b011010000_0000;
storage1[2346] = 14'b011010001_0000;
storage1[2347] = 14'b011010011_0000;
storage1[2348] = 14'b011010011_0000;
storage1[2349] = 14'b010111111_0000;
storage1[2350] = 14'b010100100_0000;
storage1[2351] = 14'b010010001_0000;
storage1[2352] = 14'b010100001_0000;
storage1[2353] = 14'b010011101_0000;
storage1[2354] = 14'b010100011_0000;
storage1[2355] = 14'b010001111_0000;
storage1[2356] = 14'b010001000_0000;
storage1[2357] = 14'b010011101_0000;
storage1[2358] = 14'b010010011_0000;
storage1[2359] = 14'b010001110_0000;
storage1[2360] = 14'b011000111_0000;
storage1[2361] = 14'b011001000_0000;
storage1[2362] = 14'b011001011_0000;
storage1[2363] = 14'b011001011_0000;
storage1[2364] = 14'b011001100_0000;
storage1[2365] = 14'b011001100_0000;
storage1[2366] = 14'b011000111_0000;
storage1[2367] = 14'b011001101_0000;
storage1[2368] = 14'b011001100_0000;
storage1[2369] = 14'b011001011_0000;
storage1[2370] = 14'b011001111_0000;
storage1[2371] = 14'b011001101_0000;
storage1[2372] = 14'b011010010_0000;
storage1[2373] = 14'b011010001_0000;
storage1[2374] = 14'b011001111_0000;
storage1[2375] = 14'b011010000_0000;
storage1[2376] = 14'b011010001_0000;
storage1[2377] = 14'b011010000_0000;
storage1[2378] = 14'b011010000_0000;
storage1[2379] = 14'b011010010_0000;
storage1[2380] = 14'b011010010_0000;
storage1[2381] = 14'b011010011_0000;
storage1[2382] = 14'b011010001_0000;
storage1[2383] = 14'b011010110_0000;
storage1[2384] = 14'b011010011_0000;
storage1[2385] = 14'b011010010_0000;
storage1[2386] = 14'b011010100_0000;
storage1[2387] = 14'b011010001_0000;
storage1[2388] = 14'b011010100_0000;
storage1[2389] = 14'b010111110_0000;
storage1[2390] = 14'b010101110_0000;
storage1[2391] = 14'b010011110_0000;
storage1[2392] = 14'b010011111_0000;
storage1[2393] = 14'b010011110_0000;
storage1[2394] = 14'b010011011_0000;
storage1[2395] = 14'b010100010_0000;
storage1[2396] = 14'b010010000_0000;
storage1[2397] = 14'b010011110_0000;
storage1[2398] = 14'b010010111_0000;
storage1[2399] = 14'b010010010_0000;
storage1[2400] = 14'b010111011_0000;
storage1[2401] = 14'b011001000_0000;
storage1[2402] = 14'b011001001_0000;
storage1[2403] = 14'b010110001_0000;
storage1[2404] = 14'b010100101_0000;
storage1[2405] = 14'b010101001_0000;
storage1[2406] = 14'b011000001_0000;
storage1[2407] = 14'b011001011_0000;
storage1[2408] = 14'b011001010_0000;
storage1[2409] = 14'b011010111_0000;
storage1[2410] = 14'b011011001_0000;
storage1[2411] = 14'b011001111_0000;
storage1[2412] = 14'b011001111_0000;
storage1[2413] = 14'b011001111_0000;
storage1[2414] = 14'b011001100_0000;
storage1[2415] = 14'b011001100_0000;
storage1[2416] = 14'b011010001_0000;
storage1[2417] = 14'b011100000_0000;
storage1[2418] = 14'b011011010_0000;
storage1[2419] = 14'b011010000_0000;
storage1[2420] = 14'b011010010_0000;
storage1[2421] = 14'b011010010_0000;
storage1[2422] = 14'b010011000_0000;
storage1[2423] = 14'b010101011_0000;
storage1[2424] = 14'b010101010_0000;
storage1[2425] = 14'b010100111_0000;
storage1[2426] = 14'b011010100_0000;
storage1[2427] = 14'b011010001_0000;
storage1[2428] = 14'b011010010_0000;
storage1[2429] = 14'b010110111_0000;
storage1[2430] = 14'b010101111_0000;
storage1[2431] = 14'b010101010_0000;
storage1[2432] = 14'b010100011_0000;
storage1[2433] = 14'b010010100_0000;
storage1[2434] = 14'b010100100_0000;
storage1[2435] = 14'b010011100_0000;
storage1[2436] = 14'b010100001_0000;
storage1[2437] = 14'b010011110_0000;
storage1[2438] = 14'b010011010_0000;
storage1[2439] = 14'b010011010_0000;
storage1[2440] = 14'b010111001_0000;
storage1[2441] = 14'b011001001_0000;
storage1[2442] = 14'b011001000_0000;
storage1[2443] = 14'b010100110_0000;
storage1[2444] = 14'b001110011_0000;
storage1[2445] = 14'b010001101_0000;
storage1[2446] = 14'b011000101_0000;
storage1[2447] = 14'b011001110_0000;
storage1[2448] = 14'b011001110_0000;
storage1[2449] = 14'b011110110_0000;
storage1[2450] = 14'b011111011_0000;
storage1[2451] = 14'b011100001_0000;
storage1[2452] = 14'b011010000_0000;
storage1[2453] = 14'b011001111_0000;
storage1[2454] = 14'b011010001_0000;
storage1[2455] = 14'b011011111_0000;
storage1[2456] = 14'b011100010_0000;
storage1[2457] = 14'b011101000_0000;
storage1[2458] = 14'b011101111_0000;
storage1[2459] = 14'b011010010_0000;
storage1[2460] = 14'b011010100_0000;
storage1[2461] = 14'b011010001_0000;
storage1[2462] = 14'b010010001_0000;
storage1[2463] = 14'b010100110_0000;
storage1[2464] = 14'b010101000_0000;
storage1[2465] = 14'b010100001_0000;
storage1[2466] = 14'b011010110_0000;
storage1[2467] = 14'b011010110_0000;
storage1[2468] = 14'b011010010_0000;
storage1[2469] = 14'b010101110_0000;
storage1[2470] = 14'b010100000_0000;
storage1[2471] = 14'b010101000_0000;
storage1[2472] = 14'b010101010_0000;
storage1[2473] = 14'b010100000_0000;
storage1[2474] = 14'b010101000_0000;
storage1[2475] = 14'b010011010_0000;
storage1[2476] = 14'b010011011_0000;
storage1[2477] = 14'b010010110_0000;
storage1[2478] = 14'b010011110_0000;
storage1[2479] = 14'b010011110_0000;
storage1[2480] = 14'b011000001_0000;
storage1[2481] = 14'b011001000_0000;
storage1[2482] = 14'b011001001_0000;
storage1[2483] = 14'b010111000_0000;
storage1[2484] = 14'b010101000_0000;
storage1[2485] = 14'b010101010_0000;
storage1[2486] = 14'b011000111_0000;
storage1[2487] = 14'b011001011_0000;
storage1[2488] = 14'b011001001_0000;
storage1[2489] = 14'b011000101_0000;
storage1[2490] = 14'b011010010_0000;
storage1[2491] = 14'b011001011_0000;
storage1[2492] = 14'b011001110_0000;
storage1[2493] = 14'b011001111_0000;
storage1[2494] = 14'b011001100_0000;
storage1[2495] = 14'b011001101_0000;
storage1[2496] = 14'b011010000_0000;
storage1[2497] = 14'b011001011_0000;
storage1[2498] = 14'b011001111_0000;
storage1[2499] = 14'b011010000_0000;
storage1[2500] = 14'b011010001_0000;
storage1[2501] = 14'b011010000_0000;
storage1[2502] = 14'b010111011_0000;
storage1[2503] = 14'b010111110_0000;
storage1[2504] = 14'b010111111_0000;
storage1[2505] = 14'b010111111_0000;
storage1[2506] = 14'b011010011_0000;
storage1[2507] = 14'b011010001_0000;
storage1[2508] = 14'b011010001_0000;
storage1[2509] = 14'b010101101_0000;
storage1[2510] = 14'b010100011_0000;
storage1[2511] = 14'b010001110_0000;
storage1[2512] = 14'b010100100_0000;
storage1[2513] = 14'b010101010_0000;
storage1[2514] = 14'b010100100_0000;
storage1[2515] = 14'b010010110_0000;
storage1[2516] = 14'b010011100_0000;
storage1[2517] = 14'b010001111_0000;
storage1[2518] = 14'b010001100_0000;
storage1[2519] = 14'b010011110_0000;
storage1[2520] = 14'b011000110_0000;
storage1[2521] = 14'b011001000_0000;
storage1[2522] = 14'b011000111_0000;
storage1[2523] = 14'b011000100_0000;
storage1[2524] = 14'b011001000_0000;
storage1[2525] = 14'b011001001_0000;
storage1[2526] = 14'b011001000_0000;
storage1[2527] = 14'b011001100_0000;
storage1[2528] = 14'b011001000_0000;
storage1[2529] = 14'b011001100_0000;
storage1[2530] = 14'b011001111_0000;
storage1[2531] = 14'b011001101_0000;
storage1[2532] = 14'b011010000_0000;
storage1[2533] = 14'b011001110_0000;
storage1[2534] = 14'b011001111_0000;
storage1[2535] = 14'b011001111_0000;
storage1[2536] = 14'b011010010_0000;
storage1[2537] = 14'b011010010_0000;
storage1[2538] = 14'b011010000_0000;
storage1[2539] = 14'b011010011_0000;
storage1[2540] = 14'b011010010_0000;
storage1[2541] = 14'b011010000_0000;
storage1[2542] = 14'b011010001_0000;
storage1[2543] = 14'b011010000_0000;
storage1[2544] = 14'b011010000_0000;
storage1[2545] = 14'b011001110_0000;
storage1[2546] = 14'b011010010_0000;
storage1[2547] = 14'b011010001_0000;
storage1[2548] = 14'b011010010_0000;
storage1[2549] = 14'b010111000_0000;
storage1[2550] = 14'b010101111_0000;
storage1[2551] = 14'b010010110_0000;
storage1[2552] = 14'b010010101_0000;
storage1[2553] = 14'b010011111_0000;
storage1[2554] = 14'b010101001_0000;
storage1[2555] = 14'b010100101_0000;
storage1[2556] = 14'b010100000_0000;
storage1[2557] = 14'b010001110_0000;
storage1[2558] = 14'b010001000_0000;
storage1[2559] = 14'b010010010_0000;
storage1[2560] = 14'b011000110_0000;
storage1[2561] = 14'b011000101_0000;
storage1[2562] = 14'b011000111_0000;
storage1[2563] = 14'b010110101_0000;
storage1[2564] = 14'b010111000_0000;
storage1[2565] = 14'b010110110_0000;
storage1[2566] = 14'b011001010_0000;
storage1[2567] = 14'b011001010_0000;
storage1[2568] = 14'b011000100_0000;
storage1[2569] = 14'b010111011_0000;
storage1[2570] = 14'b010111110_0000;
storage1[2571] = 14'b011000101_0000;
storage1[2572] = 14'b011001110_0000;
storage1[2573] = 14'b011010000_0000;
storage1[2574] = 14'b011001100_0000;
storage1[2575] = 14'b011010010_0000;
storage1[2576] = 14'b011011100_0000;
storage1[2577] = 14'b011010100_0000;
storage1[2578] = 14'b011001001_0000;
storage1[2579] = 14'b011010000_0000;
storage1[2580] = 14'b011010001_0000;
storage1[2581] = 14'b011001011_0000;
storage1[2582] = 14'b010111011_0000;
storage1[2583] = 14'b010111110_0000;
storage1[2584] = 14'b010111011_0000;
storage1[2585] = 14'b010111111_0000;
storage1[2586] = 14'b011001111_0000;
storage1[2587] = 14'b011010011_0000;
storage1[2588] = 14'b011010000_0000;
storage1[2589] = 14'b010110110_0000;
storage1[2590] = 14'b010101101_0000;
storage1[2591] = 14'b010101101_0000;
storage1[2592] = 14'b010011001_0000;
storage1[2593] = 14'b010010110_0000;
storage1[2594] = 14'b010011110_0000;
storage1[2595] = 14'b010100111_0000;
storage1[2596] = 14'b010100100_0000;
storage1[2597] = 14'b010000111_0000;
storage1[2598] = 14'b010001011_0000;
storage1[2599] = 14'b010010001_0000;
storage1[2600] = 14'b011001010_0000;
storage1[2601] = 14'b011001010_0000;
storage1[2602] = 14'b011001010_0000;
storage1[2603] = 14'b010011100_0000;
storage1[2604] = 14'b010100011_0000;
storage1[2605] = 14'b010011001_0000;
storage1[2606] = 14'b011001100_0000;
storage1[2607] = 14'b011001010_0000;
storage1[2608] = 14'b010110100_0000;
storage1[2609] = 14'b010100011_0000;
storage1[2610] = 14'b010110100_0000;
storage1[2611] = 14'b010111100_0000;
storage1[2612] = 14'b011001110_0000;
storage1[2613] = 14'b011001110_0000;
storage1[2614] = 14'b011010010_0000;
storage1[2615] = 14'b011100011_0000;
storage1[2616] = 14'b011111100_0000;
storage1[2617] = 14'b011100101_0000;
storage1[2618] = 14'b011001100_0000;
storage1[2619] = 14'b011010001_0000;
storage1[2620] = 14'b011001111_0000;
storage1[2621] = 14'b011000010_0000;
storage1[2622] = 14'b010100101_0000;
storage1[2623] = 14'b010001011_0000;
storage1[2624] = 14'b010000001_0000;
storage1[2625] = 14'b010110000_0000;
storage1[2626] = 14'b011010000_0000;
storage1[2627] = 14'b011010001_0000;
storage1[2628] = 14'b011010011_0000;
storage1[2629] = 14'b010011111_0000;
storage1[2630] = 14'b010101111_0000;
storage1[2631] = 14'b010101110_0000;
storage1[2632] = 14'b010101010_0000;
storage1[2633] = 14'b010011010_0000;
storage1[2634] = 14'b010010101_0000;
storage1[2635] = 14'b010101010_0000;
storage1[2636] = 14'b010100010_0000;
storage1[2637] = 14'b010001000_0000;
storage1[2638] = 14'b010001010_0000;
storage1[2639] = 14'b010010000_0000;
storage1[2640] = 14'b011001010_0000;
storage1[2641] = 14'b011001010_0000;
storage1[2642] = 14'b011001001_0000;
storage1[2643] = 14'b010011101_0000;
storage1[2644] = 14'b010011111_0000;
storage1[2645] = 14'b010011011_0000;
storage1[2646] = 14'b011010000_0000;
storage1[2647] = 14'b011001100_0000;
storage1[2648] = 14'b010111001_0000;
storage1[2649] = 14'b010101000_0000;
storage1[2650] = 14'b010101011_0000;
storage1[2651] = 14'b010111100_0000;
storage1[2652] = 14'b011001101_0000;
storage1[2653] = 14'b011001101_0000;
storage1[2654] = 14'b011001101_0000;
storage1[2655] = 14'b011010001_0000;
storage1[2656] = 14'b011110000_0000;
storage1[2657] = 14'b011011111_0000;
storage1[2658] = 14'b011000101_0000;
storage1[2659] = 14'b011010001_0000;
storage1[2660] = 14'b011010001_0000;
storage1[2661] = 14'b011000011_0000;
storage1[2662] = 14'b010101001_0000;
storage1[2663] = 14'b010011010_0000;
storage1[2664] = 14'b010011011_0000;
storage1[2665] = 14'b010110100_0000;
storage1[2666] = 14'b011010001_0000;
storage1[2667] = 14'b011010011_0000;
storage1[2668] = 14'b011010010_0000;
storage1[2669] = 14'b010011010_0000;
storage1[2670] = 14'b010101100_0000;
storage1[2671] = 14'b010011111_0000;
storage1[2672] = 14'b010101010_0000;
storage1[2673] = 14'b010101011_0000;
storage1[2674] = 14'b010100000_0000;
storage1[2675] = 14'b010110100_0000;
storage1[2676] = 14'b010010010_0000;
storage1[2677] = 14'b010010000_0000;
storage1[2678] = 14'b010001011_0000;
storage1[2679] = 14'b010010000_0000;
storage1[2680] = 14'b011000111_0000;
storage1[2681] = 14'b011000110_0000;
storage1[2682] = 14'b011001000_0000;
storage1[2683] = 14'b011000100_0000;
storage1[2684] = 14'b011001000_0000;
storage1[2685] = 14'b011000101_0000;
storage1[2686] = 14'b011001000_0000;
storage1[2687] = 14'b011001100_0000;
storage1[2688] = 14'b011000111_0000;
storage1[2689] = 14'b011001100_0000;
storage1[2690] = 14'b011001101_0000;
storage1[2691] = 14'b011001101_0000;
storage1[2692] = 14'b011001100_0000;
storage1[2693] = 14'b011001101_0000;
storage1[2694] = 14'b011001011_0000;
storage1[2695] = 14'b011001101_0000;
storage1[2696] = 14'b011001101_0000;
storage1[2697] = 14'b011001101_0000;
storage1[2698] = 14'b011001100_0000;
storage1[2699] = 14'b011010000_0000;
storage1[2700] = 14'b011010010_0000;
storage1[2701] = 14'b011001110_0000;
storage1[2702] = 14'b011001110_0000;
storage1[2703] = 14'b011001110_0000;
storage1[2704] = 14'b011001101_0000;
storage1[2705] = 14'b011001100_0000;
storage1[2706] = 14'b011010001_0000;
storage1[2707] = 14'b011010001_0000;
storage1[2708] = 14'b011010010_0000;
storage1[2709] = 14'b010101100_0000;
storage1[2710] = 14'b010100101_0000;
storage1[2711] = 14'b010100000_0000;
storage1[2712] = 14'b011000110_0000;
storage1[2713] = 14'b010100110_0000;
storage1[2714] = 14'b010101010_0000;
storage1[2715] = 14'b010100011_0000;
storage1[2716] = 14'b010010110_0000;
storage1[2717] = 14'b010010101_0000;
storage1[2718] = 14'b010001001_0000;
storage1[2719] = 14'b010001111_0000;
storage1[2720] = 14'b011000101_0000;
storage1[2721] = 14'b011000110_0000;
storage1[2722] = 14'b011000111_0000;
storage1[2723] = 14'b011000110_0000;
storage1[2724] = 14'b011001001_0000;
storage1[2725] = 14'b011000111_0000;
storage1[2726] = 14'b011000111_0000;
storage1[2727] = 14'b011001011_0000;
storage1[2728] = 14'b011000111_0000;
storage1[2729] = 14'b011001010_0000;
storage1[2730] = 14'b011001100_0000;
storage1[2731] = 14'b011001011_0000;
storage1[2732] = 14'b011001010_0000;
storage1[2733] = 14'b011001010_0000;
storage1[2734] = 14'b011001010_0000;
storage1[2735] = 14'b011001100_0000;
storage1[2736] = 14'b011001101_0000;
storage1[2737] = 14'b011010001_0000;
storage1[2738] = 14'b011001100_0000;
storage1[2739] = 14'b011010001_0000;
storage1[2740] = 14'b011010010_0000;
storage1[2741] = 14'b011001111_0000;
storage1[2742] = 14'b011010000_0000;
storage1[2743] = 14'b011010001_0000;
storage1[2744] = 14'b011010000_0000;
storage1[2745] = 14'b011001110_0000;
storage1[2746] = 14'b011010000_0000;
storage1[2747] = 14'b011001111_0000;
storage1[2748] = 14'b011010000_0000;
storage1[2749] = 14'b010110000_0000;
storage1[2750] = 14'b010110000_0000;
storage1[2751] = 14'b010101010_0000;
storage1[2752] = 14'b011000001_0000;
storage1[2753] = 14'b010010010_0000;
storage1[2754] = 14'b010011111_0000;
storage1[2755] = 14'b010100111_0000;
storage1[2756] = 14'b010100100_0000;
storage1[2757] = 14'b010010011_0000;
storage1[2758] = 14'b010011011_0000;
storage1[2759] = 14'b010010011_0000;
storage1[2760] = 14'b011000110_0000;
storage1[2761] = 14'b011000111_0000;
storage1[2762] = 14'b011001010_0000;
storage1[2763] = 14'b010001101_0000;
storage1[2764] = 14'b010100100_0000;
storage1[2765] = 14'b010100101_0000;
storage1[2766] = 14'b011000111_0000;
storage1[2767] = 14'b011001000_0000;
storage1[2768] = 14'b010101100_0000;
storage1[2769] = 14'b010011110_0000;
storage1[2770] = 14'b010011100_0000;
storage1[2771] = 14'b010111110_0000;
storage1[2772] = 14'b011001101_0000;
storage1[2773] = 14'b011001101_0000;
storage1[2774] = 14'b010101101_0000;
storage1[2775] = 14'b010011000_0000;
storage1[2776] = 14'b010010110_0000;
storage1[2777] = 14'b010011010_0000;
storage1[2778] = 14'b010111101_0000;
storage1[2779] = 14'b011010010_0000;
storage1[2780] = 14'b011010010_0000;
storage1[2781] = 14'b010111010_0000;
storage1[2782] = 14'b010011111_0000;
storage1[2783] = 14'b010100011_0000;
storage1[2784] = 14'b010011011_0000;
storage1[2785] = 14'b010110101_0000;
storage1[2786] = 14'b011001111_0000;
storage1[2787] = 14'b011010011_0000;
storage1[2788] = 14'b011010100_0000;
storage1[2789] = 14'b010100111_0000;
storage1[2790] = 14'b010110001_0000;
storage1[2791] = 14'b010101111_0000;
storage1[2792] = 14'b010101011_0000;
storage1[2793] = 14'b010011011_0000;
storage1[2794] = 14'b010010111_0000;
storage1[2795] = 14'b010011001_0000;
storage1[2796] = 14'b010100100_0000;
storage1[2797] = 14'b010011110_0000;
storage1[2798] = 14'b010010010_0000;
storage1[2799] = 14'b010011101_0000;
storage1[2800] = 14'b011000110_0000;
storage1[2801] = 14'b011000111_0000;
storage1[2802] = 14'b011001000_0000;
storage1[2803] = 14'b010001110_0000;
storage1[2804] = 14'b010111111_0000;
storage1[2805] = 14'b011000000_0000;
storage1[2806] = 14'b011000110_0000;
storage1[2807] = 14'b011001000_0000;
storage1[2808] = 14'b010101010_0000;
storage1[2809] = 14'b010011001_0000;
storage1[2810] = 14'b010011010_0000;
storage1[2811] = 14'b011000110_0000;
storage1[2812] = 14'b011001110_0000;
storage1[2813] = 14'b011001101_0000;
storage1[2814] = 14'b010100111_0000;
storage1[2815] = 14'b010010010_0000;
storage1[2816] = 14'b010010001_0000;
storage1[2817] = 14'b010010100_0000;
storage1[2818] = 14'b010111100_0000;
storage1[2819] = 14'b011001111_0000;
storage1[2820] = 14'b011010010_0000;
storage1[2821] = 14'b010110011_0000;
storage1[2822] = 14'b010011101_0000;
storage1[2823] = 14'b010100011_0000;
storage1[2824] = 14'b010010110_0000;
storage1[2825] = 14'b010110101_0000;
storage1[2826] = 14'b011010001_0000;
storage1[2827] = 14'b011010001_0000;
storage1[2828] = 14'b011010000_0000;
storage1[2829] = 14'b010010110_0000;
storage1[2830] = 14'b010101100_0000;
storage1[2831] = 14'b010110000_0000;
storage1[2832] = 14'b010101101_0000;
storage1[2833] = 14'b010101101_0000;
storage1[2834] = 14'b010100010_0000;
storage1[2835] = 14'b010010110_0000;
storage1[2836] = 14'b010010000_0000;
storage1[2837] = 14'b010011100_0000;
storage1[2838] = 14'b010001010_0000;
storage1[2839] = 14'b010010001_0000;
storage1[2840] = 14'b011000110_0000;
storage1[2841] = 14'b011000101_0000;
storage1[2842] = 14'b011000110_0000;
storage1[2843] = 14'b011000001_0000;
storage1[2844] = 14'b011000111_0000;
storage1[2845] = 14'b011000011_0000;
storage1[2846] = 14'b011000110_0000;
storage1[2847] = 14'b011001000_0000;
storage1[2848] = 14'b011000010_0000;
storage1[2849] = 14'b011000101_0000;
storage1[2850] = 14'b011000100_0000;
storage1[2851] = 14'b011000111_0000;
storage1[2852] = 14'b011001011_0000;
storage1[2853] = 14'b011001011_0000;
storage1[2854] = 14'b011001000_0000;
storage1[2855] = 14'b011001001_0000;
storage1[2856] = 14'b011001010_0000;
storage1[2857] = 14'b011001010_0000;
storage1[2858] = 14'b011001100_0000;
storage1[2859] = 14'b011001111_0000;
storage1[2860] = 14'b011001101_0000;
storage1[2861] = 14'b011001011_0000;
storage1[2862] = 14'b011001011_0000;
storage1[2863] = 14'b011001011_0000;
storage1[2864] = 14'b011001101_0000;
storage1[2865] = 14'b011001010_0000;
storage1[2866] = 14'b011001110_0000;
storage1[2867] = 14'b011010010_0000;
storage1[2868] = 14'b011010010_0000;
storage1[2869] = 14'b010100001_0000;
storage1[2870] = 14'b010100110_0000;
storage1[2871] = 14'b010101011_0000;
storage1[2872] = 14'b010011110_0000;
storage1[2873] = 14'b010101101_0000;
storage1[2874] = 14'b010101011_0000;
storage1[2875] = 14'b010100101_0000;
storage1[2876] = 14'b010010001_0000;
storage1[2877] = 14'b010010100_0000;
storage1[2878] = 14'b010010000_0000;
storage1[2879] = 14'b010000101_0000;
storage1[2880] = 14'b011000100_0000;
storage1[2881] = 14'b011000100_0000;
storage1[2882] = 14'b011000011_0000;
storage1[2883] = 14'b011000011_0000;
storage1[2884] = 14'b011000111_0000;
storage1[2885] = 14'b011000011_0000;
storage1[2886] = 14'b011000110_0000;
storage1[2887] = 14'b011000110_0000;
storage1[2888] = 14'b011000010_0000;
storage1[2889] = 14'b011001011_0000;
storage1[2890] = 14'b011001001_0000;
storage1[2891] = 14'b011001001_0000;
storage1[2892] = 14'b011001011_0000;
storage1[2893] = 14'b011001011_0000;
storage1[2894] = 14'b011001010_0000;
storage1[2895] = 14'b011001111_0000;
storage1[2896] = 14'b011001101_0000;
storage1[2897] = 14'b011001111_0000;
storage1[2898] = 14'b011001110_0000;
storage1[2899] = 14'b011010001_0000;
storage1[2900] = 14'b011010000_0000;
storage1[2901] = 14'b011001101_0000;
storage1[2902] = 14'b011001110_0000;
storage1[2903] = 14'b011001110_0000;
storage1[2904] = 14'b011010000_0000;
storage1[2905] = 14'b011001100_0000;
storage1[2906] = 14'b011001101_0000;
storage1[2907] = 14'b011010000_0000;
storage1[2908] = 14'b011001111_0000;
storage1[2909] = 14'b010110010_0000;
storage1[2910] = 14'b010101101_0000;
storage1[2911] = 14'b010101011_0000;
storage1[2912] = 14'b010011101_0000;
storage1[2913] = 14'b010011000_0000;
storage1[2914] = 14'b010100011_0000;
storage1[2915] = 14'b010100111_0000;
storage1[2916] = 14'b010100100_0000;
storage1[2917] = 14'b010010101_0000;
storage1[2918] = 14'b010011010_0000;
storage1[2919] = 14'b010001011_0000;
storage1[2920] = 14'b011000011_0000;
storage1[2921] = 14'b011000100_0000;
storage1[2922] = 14'b010111111_0000;
storage1[2923] = 14'b010101000_0000;
storage1[2924] = 14'b010101000_0000;
storage1[2925] = 14'b010110110_0000;
storage1[2926] = 14'b011000111_0000;
storage1[2927] = 14'b011000111_0000;
storage1[2928] = 14'b010110001_0000;
storage1[2929] = 14'b010110011_0000;
storage1[2930] = 14'b010110001_0000;
storage1[2931] = 14'b011001011_0000;
storage1[2932] = 14'b011001100_0000;
storage1[2933] = 14'b011001100_0000;
storage1[2934] = 14'b011010010_0000;
storage1[2935] = 14'b011011100_0000;
storage1[2936] = 14'b011100110_0000;
storage1[2937] = 14'b011100111_0000;
storage1[2938] = 14'b011010101_0000;
storage1[2939] = 14'b011010010_0000;
storage1[2940] = 14'b011010000_0000;
storage1[2941] = 14'b010111111_0000;
storage1[2942] = 14'b010110100_0000;
storage1[2943] = 14'b010110101_0000;
storage1[2944] = 14'b010110101_0000;
storage1[2945] = 14'b011000011_0000;
storage1[2946] = 14'b011010010_0000;
storage1[2947] = 14'b011010001_0000;
storage1[2948] = 14'b011001110_0000;
storage1[2949] = 14'b010110011_0000;
storage1[2950] = 14'b010110101_0000;
storage1[2951] = 14'b010110010_0000;
storage1[2952] = 14'b010101001_0000;
storage1[2953] = 14'b010011101_0000;
storage1[2954] = 14'b010011000_0000;
storage1[2955] = 14'b010100001_0000;
storage1[2956] = 14'b010100000_0000;
storage1[2957] = 14'b010011010_0000;
storage1[2958] = 14'b010011010_0000;
storage1[2959] = 14'b010011100_0000;
storage1[2960] = 14'b011000011_0000;
storage1[2961] = 14'b011000010_0000;
storage1[2962] = 14'b010111001_0000;
storage1[2963] = 14'b010100001_0000;
storage1[2964] = 14'b010110001_0000;
storage1[2965] = 14'b010111011_0000;
storage1[2966] = 14'b011001001_0000;
storage1[2967] = 14'b011001001_0000;
storage1[2968] = 14'b010011101_0000;
storage1[2969] = 14'b010100101_0000;
storage1[2970] = 14'b010011010_0000;
storage1[2971] = 14'b011001110_0000;
storage1[2972] = 14'b011001100_0000;
storage1[2973] = 14'b011001111_0000;
storage1[2974] = 14'b011101001_0000;
storage1[2975] = 14'b011111001_0000;
storage1[2976] = 14'b011111101_0000;
storage1[2977] = 14'b011111100_0000;
storage1[2978] = 14'b011011111_0000;
storage1[2979] = 14'b011010010_0000;
storage1[2980] = 14'b011010000_0000;
storage1[2981] = 14'b010110011_0000;
storage1[2982] = 14'b010100001_0000;
storage1[2983] = 14'b010011100_0000;
storage1[2984] = 14'b010011110_0000;
storage1[2985] = 14'b010111110_0000;
storage1[2986] = 14'b011010011_0000;
storage1[2987] = 14'b011010000_0000;
storage1[2988] = 14'b011010000_0000;
storage1[2989] = 14'b010011100_0000;
storage1[2990] = 14'b010110000_0000;
storage1[2991] = 14'b010110001_0000;
storage1[2992] = 14'b010110001_0000;
storage1[2993] = 14'b010110001_0000;
storage1[2994] = 14'b010100001_0000;
storage1[2995] = 14'b010100001_0000;
storage1[2996] = 14'b010011100_0000;
storage1[2997] = 14'b010101000_0000;
storage1[2998] = 14'b010001100_0000;
storage1[2999] = 14'b010010101_0000;
storage1[3000] = 14'b011000011_0000;
storage1[3001] = 14'b011000100_0000;
storage1[3002] = 14'b010111100_0000;
storage1[3003] = 14'b011000000_0000;
storage1[3004] = 14'b011001101_0000;
storage1[3005] = 14'b011001100_0000;
storage1[3006] = 14'b011001000_0000;
storage1[3007] = 14'b011001001_0000;
storage1[3008] = 14'b010100111_0000;
storage1[3009] = 14'b010101000_0000;
storage1[3010] = 14'b010100010_0000;
storage1[3011] = 14'b011010000_0000;
storage1[3012] = 14'b011001101_0000;
storage1[3013] = 14'b011010000_0000;
storage1[3014] = 14'b011010100_0000;
storage1[3015] = 14'b011100011_0000;
storage1[3016] = 14'b011110001_0000;
storage1[3017] = 14'b011110001_0000;
storage1[3018] = 14'b011010111_0000;
storage1[3019] = 14'b011010010_0000;
storage1[3020] = 14'b011001111_0000;
storage1[3021] = 14'b010111010_0000;
storage1[3022] = 14'b010101100_0000;
storage1[3023] = 14'b010101011_0000;
storage1[3024] = 14'b010101100_0000;
storage1[3025] = 14'b011000011_0000;
storage1[3026] = 14'b011010010_0000;
storage1[3027] = 14'b011010010_0000;
storage1[3028] = 14'b011001100_0000;
storage1[3029] = 14'b010011011_0000;
storage1[3030] = 14'b010011111_0000;
storage1[3031] = 14'b010110000_0000;
storage1[3032] = 14'b010101101_0000;
storage1[3033] = 14'b010101111_0000;
storage1[3034] = 14'b010101110_0000;
storage1[3035] = 14'b010100110_0000;
storage1[3036] = 14'b010011101_0000;
storage1[3037] = 14'b010011101_0000;
storage1[3038] = 14'b010010101_0000;
storage1[3039] = 14'b010001001_0000;
storage1[3040] = 14'b011000110_0000;
storage1[3041] = 14'b011001000_0000;
storage1[3042] = 14'b011000010_0000;
storage1[3043] = 14'b011000101_0000;
storage1[3044] = 14'b011001000_0000;
storage1[3045] = 14'b011000110_0000;
storage1[3046] = 14'b011001001_0000;
storage1[3047] = 14'b011001010_0000;
storage1[3048] = 14'b011000010_0000;
storage1[3049] = 14'b011001010_0000;
storage1[3050] = 14'b011001010_0000;
storage1[3051] = 14'b011001011_0000;
storage1[3052] = 14'b011001011_0000;
storage1[3053] = 14'b011001110_0000;
storage1[3054] = 14'b011001010_0000;
storage1[3055] = 14'b011010000_0000;
storage1[3056] = 14'b011010010_0000;
storage1[3057] = 14'b011010001_0000;
storage1[3058] = 14'b011010000_0000;
storage1[3059] = 14'b011010001_0000;
storage1[3060] = 14'b011010001_0000;
storage1[3061] = 14'b011001101_0000;
storage1[3062] = 14'b011001111_0000;
storage1[3063] = 14'b011010001_0000;
storage1[3064] = 14'b011010001_0000;
storage1[3065] = 14'b011001100_0000;
storage1[3066] = 14'b011010010_0000;
storage1[3067] = 14'b011010010_0000;
storage1[3068] = 14'b011001100_0000;
storage1[3069] = 14'b010110100_0000;
storage1[3070] = 14'b010100100_0000;
storage1[3071] = 14'b010101010_0000;
storage1[3072] = 14'b010100111_0000;
storage1[3073] = 14'b010100100_0000;
storage1[3074] = 14'b010101010_0000;
storage1[3075] = 14'b010101001_0000;
storage1[3076] = 14'b010011110_0000;
storage1[3077] = 14'b010010101_0000;
storage1[3078] = 14'b010011111_0000;
storage1[3079] = 14'b010011111_0000;
storage1[3080] = 14'b011000011_0000;
storage1[3081] = 14'b011000100_0000;
storage1[3082] = 14'b011000011_0000;
storage1[3083] = 14'b011000111_0000;
storage1[3084] = 14'b011000111_0000;
storage1[3085] = 14'b011000100_0000;
storage1[3086] = 14'b011001001_0000;
storage1[3087] = 14'b011001001_0000;
storage1[3088] = 14'b011000100_0000;
storage1[3089] = 14'b011001010_0000;
storage1[3090] = 14'b011000111_0000;
storage1[3091] = 14'b011001011_0000;
storage1[3092] = 14'b011001101_0000;
storage1[3093] = 14'b011001101_0000;
storage1[3094] = 14'b011001001_0000;
storage1[3095] = 14'b011001101_0000;
storage1[3096] = 14'b011001111_0000;
storage1[3097] = 14'b011001100_0000;
storage1[3098] = 14'b011010000_0000;
storage1[3099] = 14'b011010001_0000;
storage1[3100] = 14'b011001111_0000;
storage1[3101] = 14'b011001100_0000;
storage1[3102] = 14'b011001101_0000;
storage1[3103] = 14'b011001100_0000;
storage1[3104] = 14'b011010000_0000;
storage1[3105] = 14'b011001010_0000;
storage1[3106] = 14'b011001111_0000;
storage1[3107] = 14'b011010010_0000;
storage1[3108] = 14'b011001011_0000;
storage1[3109] = 14'b010110110_0000;
storage1[3110] = 14'b010110111_0000;
storage1[3111] = 14'b010101111_0000;
storage1[3112] = 14'b010101000_0000;
storage1[3113] = 14'b010100010_0000;
storage1[3114] = 14'b010100011_0000;
storage1[3115] = 14'b010101011_0000;
storage1[3116] = 14'b010011111_0000;
storage1[3117] = 14'b010001100_0000;
storage1[3118] = 14'b010101100_0000;
storage1[3119] = 14'b010011100_0000;
storage1[3120] = 14'b011000100_0000;
storage1[3121] = 14'b011000110_0000;
storage1[3122] = 14'b010101101_0000;
storage1[3123] = 14'b010011100_0000;
storage1[3124] = 14'b010011101_0000;
storage1[3125] = 14'b010110010_0000;
storage1[3126] = 14'b011000111_0000;
storage1[3127] = 14'b011000111_0000;
storage1[3128] = 14'b010010001_0000;
storage1[3129] = 14'b010100101_0000;
storage1[3130] = 14'b010100000_0000;
storage1[3131] = 14'b011001100_0000;
storage1[3132] = 14'b011001100_0000;
storage1[3133] = 14'b011001110_0000;
storage1[3134] = 14'b010010111_0000;
storage1[3135] = 14'b010110010_0000;
storage1[3136] = 14'b010101001_0000;
storage1[3137] = 14'b010011111_0000;
storage1[3138] = 14'b011010000_0000;
storage1[3139] = 14'b011010001_0000;
storage1[3140] = 14'b011010010_0000;
storage1[3141] = 14'b010101100_0000;
storage1[3142] = 14'b010101111_0000;
storage1[3143] = 14'b011000001_0000;
storage1[3144] = 14'b010100111_0000;
storage1[3145] = 14'b011000010_0000;
storage1[3146] = 14'b011010000_0000;
storage1[3147] = 14'b011010001_0000;
storage1[3148] = 14'b011001011_0000;
storage1[3149] = 14'b010101010_0000;
storage1[3150] = 14'b010110111_0000;
storage1[3151] = 14'b010110110_0000;
storage1[3152] = 14'b010110010_0000;
storage1[3153] = 14'b010101110_0000;
storage1[3154] = 14'b010101101_0000;
storage1[3155] = 14'b010101110_0000;
storage1[3156] = 14'b010011101_0000;
storage1[3157] = 14'b010011000_0000;
storage1[3158] = 14'b011000000_0000;
storage1[3159] = 14'b010010100_0000;
storage1[3160] = 14'b011000101_0000;
storage1[3161] = 14'b011000111_0000;
storage1[3162] = 14'b010101001_0000;
storage1[3163] = 14'b010010001_0000;
storage1[3164] = 14'b010010111_0000;
storage1[3165] = 14'b010110100_0000;
storage1[3166] = 14'b011000111_0000;
storage1[3167] = 14'b011001010_0000;
storage1[3168] = 14'b010001001_0000;
storage1[3169] = 14'b010011110_0000;
storage1[3170] = 14'b010011100_0000;
storage1[3171] = 14'b011001011_0000;
storage1[3172] = 14'b011001011_0000;
storage1[3173] = 14'b011001111_0000;
storage1[3174] = 14'b010010001_0000;
storage1[3175] = 14'b010100001_0000;
storage1[3176] = 14'b010100001_0000;
storage1[3177] = 14'b010010111_0000;
storage1[3178] = 14'b011010000_0000;
storage1[3179] = 14'b011010000_0000;
storage1[3180] = 14'b011010010_0000;
storage1[3181] = 14'b010101000_0000;
storage1[3182] = 14'b010100101_0000;
storage1[3183] = 14'b010111010_0000;
storage1[3184] = 14'b010100001_0000;
storage1[3185] = 14'b011000100_0000;
storage1[3186] = 14'b011010010_0000;
storage1[3187] = 14'b011001111_0000;
storage1[3188] = 14'b011001011_0000;
storage1[3189] = 14'b010100000_0000;
storage1[3190] = 14'b010100011_0000;
storage1[3191] = 14'b010110010_0000;
storage1[3192] = 14'b010110100_0000;
storage1[3193] = 14'b010110011_0000;
storage1[3194] = 14'b010110010_0000;
storage1[3195] = 14'b010101001_0000;
storage1[3196] = 14'b010011011_0000;
storage1[3197] = 14'b010011111_0000;
storage1[3198] = 14'b010011110_0000;
storage1[3199] = 14'b010011000_0000;

   end
   
endmodule