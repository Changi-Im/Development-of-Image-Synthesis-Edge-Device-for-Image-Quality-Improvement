module database_weight(clk,datata,re,address);

	parameter SIZE=0;

	input 							clk; 		// clock
	output	reg	signed	[SIZE-1:0]	datata;		// read data
	input 							re; 		// read signal, write signal 
	input 				[15:0] 		address;	// read address from database_weight to RAM

   
	reg signed [SIZE-1:0] storage [989:0];

	initial begin
//conv1.depthwise.depthwise.weight
storage[0] = -14'b00_00100101110;
storage[1] = 14'b00_01000101001;
storage[2] = 14'b00_01001010101;
storage[3] = 14'b00_01001110011;
storage[4] = 14'b00_01100101101;
storage[5] = -14'b00_00101110000;
storage[6] = -14'b00_01010100111;
storage[7] = 14'b00_01001111001;
storage[8] = -14'b00_00101101001;
//conv1.pointwise.pointwise.weight
storage[9] = 14'b00_00111010010;
storage[10] = -14'b01_00000100110;
storage[11] = 14'b00_11010001101;
//DB1.denseblock.0.dense_conv.depth
storage[12] = -14'b00_01000100010;
storage[13] = 14'b00_01101111001;
storage[14] = 14'b00_01000100001;
storage[15] = -14'b00_00111010000;
storage[16] = 14'b00_01011111011;
storage[17] = -14'b00_01001000001;
storage[18] = -14'b00_00011011101;
storage[19] = 14'b00_00000011001;
storage[20] = -14'b00_00010110000;
storage[21] = -14'b00_01010011101;
storage[22] = 14'b00_01000001001;
storage[23] = 14'b00_01110100101;
storage[24] = -14'b00_01010000110;
storage[25] = -14'b00_11010110000;
storage[26] = -14'b00_01111000000;
storage[27] = 14'b00_01101100111;
storage[28] = -14'b00_01010000000;
storage[29] = 14'b00_00101101100;
storage[30] = -14'b00_01010110100;
storage[31] = -14'b00_00100001100;
storage[32] = 14'b00_00110000101;
storage[33] = -14'b00_00000100011;
storage[34] = -14'b00_01000011001;
storage[35] = -14'b00_00010001000;
storage[36] = -14'b00_01100111110;
storage[37] = -14'b00_00100011110;
storage[38] = -14'b00_01001010010;
//DB1.denseblock.0.dense_conv.point
storage[39] = 14'b00_00001011111;
storage[40] = 14'b00_10010100000;
storage[41] = -14'b00_10001100101;
storage[42] = -14'b01_11010000000;
storage[43] = 14'b00_11000110101;
storage[44] = -14'b00_00011001101;
storage[45] = 14'b00_11101100101;
storage[46] = -14'b00_01011010010;
storage[47] = 14'b00_00111111010;
//DB1.denseblock.1.dense_conv.depth
storage[48] = 14'b00_01001011110;
storage[49] = 14'b00_00001001101;
storage[50] = 14'b00_00111101011;
storage[51] = 14'b00_01101000110;
storage[52] = -14'b00_00001010011;
storage[53] = 14'b00_00001000101;
storage[54] = -14'b00_00010101011;
storage[55] = 14'b00_00101111000;
storage[56] = 14'b00_00110100111;
storage[57] = -14'b00_00010110011;
storage[58] = 14'b00_00010010001;
storage[59] = 14'b01_01101010110;
storage[60] = -14'b00_00001100001;
storage[61] = 14'b00_00110101101;
storage[62] = 14'b00_00001001000;
storage[63] = 14'b00_11000111110;
storage[64] = 14'b00_10110111010;
storage[65] = 14'b00_11000010000;
storage[66] = 14'b00_01010000111;
storage[67] = 14'b00_10010111001;
storage[68] = -14'b00_00000111001;
storage[69] = 14'b00_10001110010;
storage[70] = 14'b00_00001001111;
storage[71] = -14'b00_00101111101;
storage[72] = 14'b00_00100110001;
storage[73] = 14'b00_01001100010;
storage[74] = 14'b00_00011001101;
storage[75] = 14'b00_01001010010;
storage[76] = 14'b00_00000101101;
storage[77] = -14'b00_00101010101;
storage[78] = 14'b00_01010100110;
storage[79] = 14'b00_00100011000;
storage[80] = 14'b00_00000010010;
storage[81] = 14'b00_00111110110;
storage[82] = 14'b00_00001110111;
storage[83] = 14'b00_01011101010;
storage[84] = -14'b00_00110101011;
storage[85] = -14'b00_00111110100;
storage[86] = -14'b00_00101101111;
storage[87] = -14'b00_01011010110;
storage[88] = 14'b00_00011100101;
storage[89] = -14'b00_01111001010;
storage[90] = 14'b00_00011111011;
storage[91] = -14'b00_00010001110;
storage[92] = -14'b00_01000000101;
storage[93] = 14'b00_01000110011;
storage[94] = 14'b00_00001111111;
storage[95] = 14'b01_00000010110;
storage[96] = -14'b00_00000111001;
storage[97] = 14'b00_00011100000;
storage[98] = 14'b00_10110110011;
storage[99] = 14'b00_00110011011;
storage[100] = 14'b00_01100101011;
storage[101] = 14'b00_11110010101;
//DB1.denseblock.1.dense_conv.point
storage[102] = -14'b00_00001101010;
storage[103] = 14'b00_10010011111;
storage[104] = 14'b00_00111011111;
storage[105] = 14'b00_00110011001;
storage[106] = -14'b00_10010001001;
storage[107] = 14'b00_10011011111;
storage[108] = 14'b00_01111001111;
storage[109] = -14'b10_00010100000;
storage[110] = 14'b00_01011111111;
storage[111] = 14'b00_01011101011;
storage[112] = 14'b00_00110011101;
storage[113] = -14'b00_01010010100;
storage[114] = 14'b00_00011011000;
storage[115] = -14'b00_01000110010;
storage[116] = 14'b00_01101011001;
storage[117] = -14'b00_00000110000;
storage[118] = -14'b00_01110000110;
storage[119] = -14'b01_01000100000;
//DB1.denseblock.2.dense_conv.depth
storage[120] = -14'b00_11111010100;
storage[121] = -14'b00_00011111000;
storage[122] = 14'b00_11010110011;
storage[123] = 14'b00_00111001110;
storage[124] = -14'b00_00001010101;
storage[125] = 14'b00_01011011001;
storage[126] = -14'b00_11001100101;
storage[127] = -14'b01_00111001100;
storage[128] = -14'b00_00010100011;
storage[129] = 14'b00_01111110010;
storage[130] = 14'b00_01110111010;
storage[131] = -14'b00_00000011111;
storage[132] = 14'b00_11000110101;
storage[133] = -14'b00_00101100101;
storage[134] = -14'b00_10110000001;
storage[135] = 14'b00_01111110001;
storage[136] = -14'b00_01100100010;
storage[137] = -14'b00_00110110100;
storage[138] = 14'b00_00011100100;
storage[139] = 14'b00_01000110100;
storage[140] = -14'b00_00111001111;
storage[141] = 14'b00_01000010001;
storage[142] = -14'b00_01000001111;
storage[143] = -14'b00_01001000011;
storage[144] = 14'b00_00011110010;
storage[145] = -14'b00_00110110111;
storage[146] = -14'b00_01110101101;
storage[147] = -14'b00_00111010111;
storage[148] = 14'b00_00111011100;
storage[149] = 14'b00_00010101011;
storage[150] = -14'b00_00111111100;
storage[151] = 14'b00_01100000101;
storage[152] = 14'b00_01100110111;
storage[153] = 14'b00_00100000000;
storage[154] = 14'b00_00100010001;
storage[155] = 14'b00_00010101011;
storage[156] = 14'b00_01100100111;
storage[157] = -14'b00_01100010011;
storage[158] = -14'b00_00100001000;
storage[159] = -14'b00_10001110111;
storage[160] = -14'b00_01000101000;
storage[161] = -14'b00_01110100111;
storage[162] = -14'b00_11010000111;
storage[163] = 14'b00_00110111100;
storage[164] = -14'b00_01100011101;
storage[165] = -14'b00_11110110110;
storage[166] = -14'b00_10000111100;
storage[167] = -14'b00_10100100111;
storage[168] = -14'b01_00000110100;
storage[169] = -14'b00_10101101110;
storage[170] = -14'b00_11011000010;
storage[171] = -14'b00_10100000111;
storage[172] = -14'b01_00111101000;
storage[173] = -14'b01_01001001010;
storage[174] = 14'b00_00111011000;
storage[175] = -14'b00_00111000001;
storage[176] = 14'b00_01001001100;
storage[177] = 14'b00_00001010010;
storage[178] = -14'b00_00000111110;
storage[179] = -14'b00_01011010010;
storage[180] = 14'b00_00100100100;
storage[181] = 14'b00_00100111010;
storage[182] = 14'b00_00111000010;
storage[183] = -14'b00_00111111111;
storage[184] = 14'b00_00101110000;
storage[185] = -14'b00_00011011010;
storage[186] = -14'b00_00001011001;
storage[187] = 14'b00_00000001000;
storage[188] = -14'b00_00000000010;
storage[189] = -14'b00_00110101000;
storage[190] = 14'b00_00100001110;
storage[191] = -14'b00_01010100011;
storage[192] = 14'b00_00001100110;
storage[193] = 14'b00_00101111100;
storage[194] = 14'b00_00110100100;
storage[195] = -14'b00_00110001100;
storage[196] = 14'b00_00010001001;
storage[197] = 14'b00_01010010010;
storage[198] = -14'b00_00000101111;
storage[199] = -14'b00_00110101100;
storage[200] = 14'b00_00111010000;
//DB1.denseblock.2.dense_conv.point
storage[201] = -14'b00_01101110001;
storage[202] = 14'b00_11000000000;
storage[203] = -14'b00_10010010000;
storage[204] = 14'b00_00100011000;
storage[205] = -14'b00_01010010010;
storage[206] = -14'b00_00111100001;
storage[207] = -14'b00_00110000000;
storage[208] = -14'b00_00010000000;
storage[209] = 14'b00_00010010101;
storage[210] = -14'b00_01001110101;
storage[211] = -14'b00_00101111010;
storage[212] = 14'b00_00010111011;
storage[213] = 14'b00_00000010100;
storage[214] = -14'b00_00101011110;
storage[215] = 14'b01_00010001010;
storage[216] = 14'b00_01000000011;
storage[217] = -14'b00_01000000100;
storage[218] = -14'b00_00001010010;
storage[219] = 14'b00_00000111110;
storage[220] = 14'b00_00011000000;
storage[221] = -14'b00_00101110100;
storage[222] = 14'b00_00010111110;
storage[223] = 14'b00_00010010011;
storage[224] = 14'b00_10001110110;
storage[225] = -14'b00_01110000010;
storage[226] = -14'b00_01011110101;
storage[227] = -14'b00_11100100110;
//conv1_1.depthwise.depthwise.weigh
storage[228] = 14'b00_01001110110;
storage[229] = -14'b00_00110010101;
storage[230] = -14'b00_00100110100;
storage[231] = 14'b00_01010111101;
storage[232] = 14'b00_01101111011;
storage[233] = -14'b00_00101011000;
storage[234] = 14'b00_01010111100;
storage[235] = 14'b00_00101000011;
storage[236] = 14'b00_00111010101;
//conv1_1.pointwise.pointwise.weigh
storage[237] = 14'b00_01101000100;
storage[238] = 14'b00_01111010010;
storage[239] = -14'b01_01010001010;
//DB2.denseblock.0.dense_conv.depth
storage[240] = 14'b00_01001110001;
storage[241] = -14'b00_00011000000;
storage[242] = 14'b00_00011011010;
storage[243] = 14'b00_00011100101;
storage[244] = -14'b00_00010110011;
storage[245] = 14'b00_00110101111;
storage[246] = -14'b00_00000111110;
storage[247] = 14'b00_01100110100;
storage[248] = 14'b00_00101011001;
storage[249] = 14'b00_00000110011;
storage[250] = -14'b00_00111011111;
storage[251] = 14'b00_01110001111;
storage[252] = -14'b00_00110010111;
storage[253] = -14'b00_01011001000;
storage[254] = -14'b00_01001110011;
storage[255] = -14'b00_01100011000;
storage[256] = 14'b00_00110010101;
storage[257] = -14'b00_00100001100;
storage[258] = -14'b00_10001010111;
storage[259] = -14'b00_01101101110;
storage[260] = 14'b00_00111010000;
storage[261] = -14'b00_11000100011;
storage[262] = 14'b00_00001000100;
storage[263] = -14'b00_01110001010;
storage[264] = -14'b01_00001010100;
storage[265] = -14'b00_00111101001;
storage[266] = -14'b00_01011011101;
//DB2.denseblock.0.dense_conv.point
storage[267] = 14'b00_01101001001;
storage[268] = 14'b00_01101000111;
storage[269] = 14'b00_11011011010;
storage[270] = 14'b00_01001110111;
storage[271] = -14'b00_01101111010;
storage[272] = -14'b00_00101001011;
storage[273] = -14'b00_00111000011;
storage[274] = -14'b00_10001001010;
storage[275] = 14'b00_00000111001;
//DB2.denseblock.1.dense_conv.depth
storage[276] = 14'b00_01110011111;
storage[277] = -14'b00_00100001011;
storage[278] = 14'b00_01100110100;
storage[279] = 14'b00_01101010111;
storage[280] = 14'b00_00110011001;
storage[281] = -14'b00_00100101001;
storage[282] = -14'b00_00011000110;
storage[283] = 14'b00_01000111101;
storage[284] = 14'b00_01000011010;
storage[285] = 14'b00_00101001100;
storage[286] = -14'b00_01000001001;
storage[287] = -14'b00_00011101101;
storage[288] = 14'b00_00110000100;
storage[289] = -14'b00_00101101110;
storage[290] = 14'b00_01110110001;
storage[291] = -14'b00_00010111010;
storage[292] = -14'b00_00101001110;
storage[293] = 14'b00_01010111100;
storage[294] = -14'b01_00010001000;
storage[295] = -14'b00_01101001100;
storage[296] = 14'b00_00110000100;
storage[297] = 14'b00_00110001111;
storage[298] = -14'b00_01011100000;
storage[299] = 14'b00_01111100000;
storage[300] = 14'b00_01001100000;
storage[301] = 14'b00_10000010110;
storage[302] = -14'b00_01010001101;
storage[303] = -14'b00_00010011110;
storage[304] = 14'b01_00101001110;
storage[305] = 14'b00_11000010001;
storage[306] = -14'b00_10101000101;
storage[307] = 14'b00_10011111001;
storage[308] = 14'b00_01001111110;
storage[309] = -14'b00_00100100000;
storage[310] = 14'b01_01101100110;
storage[311] = 14'b00_11111111100;
storage[312] = -14'b00_00011100011;
storage[313] = 14'b00_00010101110;
storage[314] = -14'b00_00100111000;
storage[315] = 14'b00_00001110110;
storage[316] = -14'b00_01001100111;
storage[317] = 14'b00_00111110100;
storage[318] = 14'b00_00101001100;
storage[319] = -14'b00_00011110100;
storage[320] = -14'b00_00111011001;
storage[321] = 14'b00_00110100000;
storage[322] = 14'b00_00101101001;
storage[323] = 14'b00_00100011001;
storage[324] = 14'b00_00011111100;
storage[325] = 14'b00_00010010010;
storage[326] = 14'b00_00111011000;
storage[327] = 14'b00_00001010001;
storage[328] = -14'b00_00000101101;
storage[329] = -14'b00_00101101011;
//DB2.denseblock.1.dense_conv.point
storage[330] = -14'b00_00010101010;
storage[331] = 14'b00_01011110000;
storage[332] = 14'b00_01100100011;
storage[333] = -14'b00_00000111110;
storage[334] = -14'b00_01000111011;
storage[335] = -14'b00_00011011100;
storage[336] = 14'b00_01000000011;
storage[337] = 14'b00_00100111100;
storage[338] = -14'b00_10110010010;
storage[339] = 14'b01_00110111000;
storage[340] = 14'b00_01100011110;
storage[341] = -14'b00_00000010101;
storage[342] = 14'b00_01001011000;
storage[343] = 14'b00_00111111111;
storage[344] = 14'b00_01101111001;
storage[345] = 14'b10_01000101100;
storage[346] = -14'b00_01101111001;
storage[347] = 14'b00_00100100111;
//DB2.denseblock.2.dense_conv.depth
storage[348] = 14'b00_00011111101;
storage[349] = 14'b00_01001011100;
storage[350] = 14'b00_01011011001;
storage[351] = -14'b00_00111111110;
storage[352] = -14'b00_00101000000;
storage[353] = 14'b00_00100111111;
storage[354] = 14'b00_00101010010;
storage[355] = -14'b00_00100110001;
storage[356] = 14'b00_00000000110;
storage[357] = -14'b00_00111010011;
storage[358] = -14'b00_00011101100;
storage[359] = -14'b00_00001001100;
storage[360] = -14'b00_00011010111;
storage[361] = 14'b00_00011010101;
storage[362] = 14'b00_00001010000;
storage[363] = -14'b00_01000000001;
storage[364] = -14'b00_00111101111;
storage[365] = -14'b00_01010010101;
storage[366] = 14'b00_00110000010;
storage[367] = 14'b00_10101100101;
storage[368] = 14'b00_10011101011;
storage[369] = 14'b00_00011111000;
storage[370] = -14'b00_00001101010;
storage[371] = 14'b00_01110110000;
storage[372] = -14'b00_01010001010;
storage[373] = -14'b00_11100111010;
storage[374] = 14'b00_00010001101;
storage[375] = -14'b00_11000011010;
storage[376] = 14'b00_01001000011;
storage[377] = -14'b00_10001111111;
storage[378] = -14'b00_01110011011;
storage[379] = 14'b00_01110101000;
storage[380] = -14'b00_10110010111;
storage[381] = -14'b00_00101010101;
storage[382] = 14'b00_01001101000;
storage[383] = -14'b00_01110001000;
storage[384] = -14'b00_00001011111;
storage[385] = 14'b00_00110110001;
storage[386] = 14'b00_00010000100;
storage[387] = -14'b00_01001011101;
storage[388] = -14'b00_00100111000;
storage[389] = 14'b00_00001111011;
storage[390] = -14'b00_00100100001;
storage[391] = 14'b00_01000001001;
storage[392] = -14'b00_01010100110;
storage[393] = 14'b00_00101101011;
storage[394] = -14'b00_00011101100;
storage[395] = 14'b00_01000111110;
storage[396] = -14'b00_00111110010;
storage[397] = -14'b00_00010100010;
storage[398] = -14'b00_01000001101;
storage[399] = 14'b00_01000110010;
storage[400] = 14'b00_00110000111;
storage[401] = -14'b00_00010101000;
storage[402] = -14'b00_01101111001;
storage[403] = -14'b00_10000011110;
storage[404] = 14'b00_01001000110;
storage[405] = -14'b00_00000100000;
storage[406] = -14'b00_11101001011;
storage[407] = 14'b00_01111110000;
storage[408] = 14'b00_01100111110;
storage[409] = -14'b00_00101101100;
storage[410] = 14'b00_10111110101;
storage[411] = 14'b00_01010110011;
storage[412] = -14'b00_00001010111;
storage[413] = 14'b00_01010111010;
storage[414] = -14'b00_00001010010;
storage[415] = 14'b00_00001111010;
storage[416] = 14'b00_01001111011;
storage[417] = 14'b00_00001010101;
storage[418] = -14'b00_00100001101;
storage[419] = 14'b00_00100011010;
storage[420] = -14'b00_01001100011;
storage[421] = -14'b00_00110101010;
storage[422] = 14'b00_00101101111;
storage[423] = 14'b00_00011110001;
storage[424] = 14'b00_00110101110;
storage[425] = 14'b00_01010001100;
storage[426] = -14'b00_00000100101;
storage[427] = -14'b00_00110011110;
storage[428] = -14'b00_00011010100;
//DB2.denseblock.2.dense_conv.point
storage[429] = 14'b00_01010011001;
storage[430] = -14'b00_00001000100;
storage[431] = -14'b00_10101010100;
storage[432] = 14'b00_10101101111;
storage[433] = 14'b00_00101010000;
storage[434] = -14'b00_00010110000;
storage[435] = -14'b00_11111101010;
storage[436] = 14'b00_00011111110;
storage[437] = 14'b00_11000001000;
storage[438] = -14'b00_00010010000;
storage[439] = -14'b00_00011001101;
storage[440] = 14'b01_00011000010;
storage[441] = -14'b01_00000000110;
storage[442] = -14'b00_00110000000;
storage[443] = 14'b00_00010000011;
storage[444] = 14'b00_01111010000;
storage[445] = 14'b00_01001100001;
storage[446] = -14'b00_00001001000;
storage[447] = -14'b00_00100000011;
storage[448] = -14'b00_00101010100;
storage[449] = 14'b01_10101000110;
storage[450] = -14'b00_01101110101;
storage[451] = -14'b00_00100110011;
storage[452] = 14'b00_00110101011;
storage[453] = -14'b00_11001100010;
storage[454] = 14'b00_00110101101;
storage[455] = 14'b00_11010100101;
//conv2.depthwise.depthwise.weight
storage[456] = -14'b00_00011100110;
storage[457] = 14'b00_01101001100;
storage[458] = 14'b00_01011001001;
storage[459] = 14'b00_01011001011;
storage[460] = -14'b00_00001101010;
storage[461] = 14'b00_00010001110;
storage[462] = 14'b00_00111000111;
storage[463] = -14'b00_00000111011;
storage[464] = 14'b00_00101000011;
storage[465] = -14'b00_00100101011;
storage[466] = 14'b00_00111001011;
storage[467] = 14'b00_01000101111;
storage[468] = -14'b00_00010011111;
storage[469] = -14'b00_00111111100;
storage[470] = 14'b00_01101001000;
storage[471] = -14'b00_00001011110;
storage[472] = -14'b00_00010101111;
storage[473] = -14'b00_00100011111;
storage[474] = -14'b00_01000111110;
storage[475] = -14'b00_01101111001;
storage[476] = -14'b00_01000010100;
storage[477] = -14'b00_01001110111;
storage[478] = 14'b01_01000100100;
storage[479] = -14'b00_00110101011;
storage[480] = -14'b00_00001111101;
storage[481] = -14'b01_00010111010;
storage[482] = 14'b00_00101011011;
storage[483] = -14'b00_00011101111;
storage[484] = -14'b00_00001110101;
storage[485] = -14'b00_01000001010;
storage[486] = -14'b00_00010101010;
storage[487] = -14'b00_01010100001;
storage[488] = -14'b00_01001000110;
storage[489] = -14'b00_00011100100;
storage[490] = 14'b00_00010101111;
storage[491] = 14'b00_00100101001;
storage[492] = 14'b00_01000011100;
storage[493] = -14'b00_01001101101;
storage[494] = 14'b00_01010011100;
storage[495] = 14'b00_00011110100;
storage[496] = 14'b00_00011110011;
storage[497] = -14'b00_00011110110;
storage[498] = -14'b00_01011111010;
storage[499] = -14'b00_00011000110;
storage[500] = -14'b00_00010111001;
storage[501] = -14'b00_01000001100;
storage[502] = -14'b00_00001110111;
storage[503] = -14'b00_01001111111;
storage[504] = 14'b00_00101101011;
storage[505] = -14'b00_00010111111;
storage[506] = -14'b00_00001000100;
storage[507] = 14'b00_00110001001;
storage[508] = 14'b00_00011100001;
storage[509] = 14'b00_00101010101;
storage[510] = -14'b00_00010010011;
storage[511] = -14'b00_01100100010;
storage[512] = -14'b00_00110001010;
storage[513] = 14'b00_00011000000;
storage[514] = -14'b00_00101011110;
storage[515] = -14'b00_01010001110;
storage[516] = 14'b00_00101000101;
storage[517] = -14'b00_01010000001;
storage[518] = 14'b00_01000100100;
storage[519] = -14'b00_00001110100;
storage[520] = -14'b00_00100011110;
storage[521] = -14'b00_10010001010;
storage[522] = 14'b00_01011011111;
storage[523] = 14'b00_01110111010;
storage[524] = -14'b00_00100101110;
storage[525] = 14'b00_00001010110;
storage[526] = -14'b00_00010000101;
storage[527] = 14'b00_00101100111;
storage[528] = -14'b00_00011101011;
storage[529] = -14'b00_01101101111;
storage[530] = -14'b00_10001011101;
storage[531] = -14'b00_01000011010;
storage[532] = 14'b00_00010111000;
storage[533] = -14'b00_01010110111;
storage[534] = 14'b00_00000001010;
storage[535] = 14'b00_00001001000;
storage[536] = -14'b00_01001101000;
storage[537] = -14'b00_00101000010;
storage[538] = -14'b00_01111100011;
storage[539] = 14'b00_00000011001;
storage[540] = -14'b00_00101011100;
storage[541] = -14'b00_00110001101;
storage[542] = 14'b00_00110100100;
storage[543] = -14'b00_00000101101;
storage[544] = 14'b00_00010101110;
storage[545] = 14'b00_00100001010;
storage[546] = 14'b00_00101101100;
storage[547] = 14'b00_00011000011;
storage[548] = 14'b00_00010111000;
storage[549] = 14'b00_00100100101;
storage[550] = 14'b00_01000110010;
storage[551] = -14'b00_00110111010;
storage[552] = 14'b00_01110110000;
storage[553] = 14'b00_00111110000;
storage[554] = -14'b00_00000110110;
storage[555] = -14'b00_00110110100;
storage[556] = 14'b00_00101001100;
storage[557] = 14'b00_00110100000;
storage[558] = -14'b00_01000101001;
storage[559] = -14'b00_00010101101;
storage[560] = -14'b00_00111010011;
storage[561] = -14'b00_00010000111;
storage[562] = -14'b00_00100111010;
storage[563] = 14'b00_00000000110;
//conv2.pointwise.pointwise.weight
storage[564] = 14'b00_00100001100;
storage[565] = -14'b00_10000010101;
storage[566] = 14'b00_00101100010;
storage[567] = -14'b00_01010100101;
storage[568] = 14'b00_00000101001;
storage[569] = -14'b00_00001111100;
storage[570] = -14'b00_01001001101;
storage[571] = 14'b00_10101111110;
storage[572] = 14'b00_01010001101;
storage[573] = -14'b00_00000100001;
storage[574] = -14'b00_10100000111;
storage[575] = -14'b00_01010010100;
storage[576] = -14'b00_00000000000;
storage[577] = -14'b00_00011110000;
storage[578] = 14'b00_00010110011;
storage[579] = 14'b00_01001100101;
storage[580] = -14'b00_00011001111;
storage[581] = 14'b00_00101011001;
storage[582] = -14'b00_00001010001;
storage[583] = -14'b00_00100110101;
storage[584] = -14'b00_00001100110;
storage[585] = 14'b00_00001111110;
storage[586] = 14'b00_00010001001;
storage[587] = -14'b00_01001100101;
storage[588] = 14'b00_01000001110;
storage[589] = 14'b00_01001111100;
storage[590] = 14'b00_00000100010;
storage[591] = -14'b00_01000100110;
storage[592] = 14'b00_00101011001;
storage[593] = -14'b00_00010000010;
storage[594] = -14'b00_00000101110;
storage[595] = -14'b00_00100101000;
storage[596] = -14'b00_00010101110;
storage[597] = -14'b00_01000111011;
storage[598] = -14'b00_00111011001;
storage[599] = 14'b00_00011111101;
storage[600] = 14'b00_00010100111;
storage[601] = 14'b00_01010100000;
storage[602] = -14'b00_01000000011;
storage[603] = -14'b00_00111000110;
storage[604] = 14'b00_00110000100;
storage[605] = -14'b00_01111110000;
storage[606] = -14'b00_00111001110;
storage[607] = 14'b00_00100111011;
storage[608] = -14'b00_01001000010;
storage[609] = 14'b00_00110111110;
storage[610] = -14'b00_00110100001;
storage[611] = -14'b00_00100001111;
storage[612] = 14'b00_01010110001;
storage[613] = -14'b00_00110011100;
storage[614] = 14'b00_00000010111;
storage[615] = -14'b00_00001111010;
storage[616] = 14'b00_00001010111;
storage[617] = -14'b00_01101010111;
storage[618] = -14'b00_00111001100;
storage[619] = 14'b00_00010000101;
storage[620] = 14'b00_00101011111;
storage[621] = -14'b00_01000011001;
storage[622] = -14'b00_01100010001;
storage[623] = 14'b00_01001000000;
storage[624] = -14'b00_00100001111;
storage[625] = -14'b00_01001101101;
storage[626] = -14'b00_00001110001;
storage[627] = -14'b00_00100010010;
storage[628] = 14'b00_00010100001;
storage[629] = 14'b00_00100011011;
storage[630] = -14'b00_00001101100;
storage[631] = -14'b00_00101000001;
storage[632] = -14'b00_01010000101;
storage[633] = 14'b00_10000110000;
storage[634] = 14'b00_00000101000;
storage[635] = -14'b00_00101010110;
storage[636] = -14'b00_00000011100;
storage[637] = 14'b00_01010010000;
storage[638] = 14'b00_00000010100;
storage[639] = -14'b00_00011010011;
storage[640] = -14'b00_00011101000;
storage[641] = 14'b00_00010000000;
storage[642] = -14'b00_00101100001;
storage[643] = -14'b00_00001111010;
storage[644] = -14'b00_00011000101;
storage[645] = -14'b00_01001100101;
storage[646] = -14'b00_00010011000;
storage[647] = 14'b00_00011111110;
storage[648] = 14'b00_10111011111;
storage[649] = 14'b10_01010110100;
storage[650] = 14'b10_00101111100;
storage[651] = -14'b01_00010101110;
storage[652] = -14'b10_00100110000;
storage[653] = -14'b01_00011100000;
storage[654] = -14'b01_00011100000;
storage[655] = -14'b00_10110010011;
storage[656] = -14'b00_00010010010;
storage[657] = -14'b01_10101000110;
storage[658] = 14'b00_00111101011;
storage[659] = 14'b00_11011111000;
storage[660] = 14'b00_00110101000;
storage[661] = 14'b00_00101011101;
storage[662] = -14'b00_00111110111;
storage[663] = -14'b00_01000000110;
storage[664] = 14'b00_00111011111;
storage[665] = -14'b00_00010010100;
storage[666] = -14'b00_01000111100;
storage[667] = -14'b00_00000000101;
storage[668] = -14'b00_01010010100;
storage[669] = -14'b00_01010101100;
storage[670] = 14'b00_00010110100;
storage[671] = 14'b00_00100111111;
storage[672] = 14'b00_01000011101;
storage[673] = 14'b00_01001101101;
storage[674] = -14'b00_00100010001;
storage[675] = -14'b00_01000111110;
storage[676] = 14'b00_00000001000;
storage[677] = -14'b00_01011000010;
storage[678] = -14'b00_00101101110;
storage[679] = 14'b00_00111111011;
storage[680] = 14'b00_00110011011;
storage[681] = -14'b00_00110110110;
storage[682] = -14'b00_00010110101;
storage[683] = 14'b00_00000110000;
storage[684] = 14'b00_01010011101;
storage[685] = 14'b00_01010100000;
storage[686] = 14'b00_00011100101;
storage[687] = -14'b00_00111101100;
storage[688] = -14'b00_00100111011;
storage[689] = -14'b00_00010111001;
storage[690] = -14'b00_01011101011;
storage[691] = -14'b00_00001110110;
storage[692] = 14'b00_00100110110;
storage[693] = -14'b00_00101111111;
storage[694] = -14'b00_01101101110;
storage[695] = 14'b00_00001000011;
storage[696] = 14'b00_00100110010;
storage[697] = 14'b00_00101001111;
storage[698] = -14'b00_00100100000;
storage[699] = -14'b00_00001111001;
storage[700] = 14'b00_01000011011;
storage[701] = -14'b00_00011100000;
storage[702] = 14'b00_00000011000;
storage[703] = 14'b00_01000111110;
storage[704] = -14'b00_01010010011;
storage[705] = -14'b00_00001011010;
storage[706] = -14'b00_00111010100;
storage[707] = 14'b00_01000101100;
//conv3.depthwise.depthwise.weight
storage[708] = 14'b00_00010111101;
storage[709] = 14'b01_11011001000;
storage[710] = 14'b00_10001110101;
storage[711] = 14'b01_10100011000;
storage[712] = 14'b10_00011101000;
storage[713] = 14'b00_00111111000;
storage[714] = 14'b00_01010111110;
storage[715] = 14'b01_00110010000;
storage[716] = -14'b01_10000101100;
storage[717] = -14'b00_00101110100;
storage[718] = 14'b00_00000001000;
storage[719] = -14'b00_10001000111;
storage[720] = -14'b00_01100101011;
storage[721] = -14'b00_10001110011;
storage[722] = -14'b00_00111100000;
storage[723] = -14'b00_01100101000;
storage[724] = -14'b00_00010010111;
storage[725] = -14'b00_00000011001;
storage[726] = -14'b00_01110110010;
storage[727] = -14'b00_00011101010;
storage[728] = -14'b00_00101011100;
storage[729] = -14'b00_01001101000;
storage[730] = -14'b00_01101111101;
storage[731] = -14'b00_00101010100;
storage[732] = -14'b00_00110110001;
storage[733] = -14'b00_00100101111;
storage[734] = 14'b00_00010111000;
storage[735] = 14'b00_00000111010;
storage[736] = -14'b00_01011000011;
storage[737] = 14'b00_00001111101;
storage[738] = 14'b00_00100001001;
storage[739] = -14'b00_00011001111;
storage[740] = 14'b00_00001001100;
storage[741] = -14'b00_00101001110;
storage[742] = 14'b00_00001001011;
storage[743] = -14'b00_01011011000;
storage[744] = -14'b00_00110111010;
storage[745] = 14'b00_00011100101;
storage[746] = -14'b00_01110000100;
storage[747] = -14'b00_00111000111;
storage[748] = -14'b00_00100010110;
storage[749] = -14'b00_00011010001;
storage[750] = -14'b00_00011011101;
storage[751] = 14'b00_00010110101;
storage[752] = -14'b00_01001011001;
storage[753] = -14'b00_00110000100;
storage[754] = 14'b00_10000010011;
storage[755] = 14'b00_01010110010;
storage[756] = 14'b00_01000011001;
storage[757] = 14'b00_01110010100;
storage[758] = -14'b00_00010010100;
storage[759] = 14'b00_10000110001;
storage[760] = 14'b00_00000100001;
storage[761] = -14'b00_01101110111;
storage[762] = 14'b00_00010010001;
storage[763] = 14'b00_00100010001;
storage[764] = -14'b00_01000110111;
storage[765] = 14'b00_00001110010;
storage[766] = 14'b00_01000010010;
storage[767] = -14'b00_00111110000;
storage[768] = 14'b00_01111001000;
storage[769] = 14'b00_01111110010;
storage[770] = 14'b00_00111100001;
storage[771] = -14'b00_00000101101;
storage[772] = -14'b00_01101000100;
storage[773] = 14'b00_01001011000;
storage[774] = -14'b00_00001000000;
storage[775] = -14'b00_10010111000;
storage[776] = -14'b00_10000110010;
storage[777] = 14'b00_10000100100;
storage[778] = 14'b00_00001100011;
storage[779] = 14'b00_10101010010;
storage[780] = 14'b00_00011100000;
storage[781] = -14'b00_01101000011;
storage[782] = 14'b00_00000100001;
storage[783] = -14'b00_00110111000;
storage[784] = 14'b00_00000101001;
storage[785] = -14'b00_00000110010;
storage[786] = -14'b00_00000001000;
storage[787] = -14'b00_01001111110;
storage[788] = -14'b00_01001110111;
storage[789] = -14'b00_00001100100;
storage[790] = 14'b00_00100101110;
storage[791] = 14'b00_01110001101;
storage[792] = 14'b00_01000110011;
storage[793] = 14'b00_01000011110;
storage[794] = -14'b00_00001000001;
storage[795] = -14'b00_00001101101;
storage[796] = -14'b00_00010011111;
storage[797] = 14'b00_01011101011;
storage[798] = 14'b00_00000001011;
storage[799] = -14'b00_01011100110;
storage[800] = 14'b00_00100111011;
storage[801] = -14'b00_00000000110;
storage[802] = 14'b00_00001111100;
storage[803] = -14'b00_01110100110;
storage[804] = -14'b00_01101110000;
storage[805] = -14'b00_01101000100;
storage[806] = -14'b00_01010110100;
storage[807] = -14'b00_01001110110;
storage[808] = -14'b00_00100000011;
storage[809] = -14'b00_01011111001;
storage[810] = 14'b00_00001110100;
storage[811] = -14'b00_01000101100;
storage[812] = -14'b00_01100100110;
storage[813] = -14'b00_00111101011;
storage[814] = -14'b00_01010110101;
storage[815] = -14'b00_01010100100;
//conv3.pointwise.pointwise.weight
storage[816] = 14'b00_10100011010;
storage[817] = -14'b00_01000111110;
storage[818] = 14'b00_00001111010;
storage[819] = 14'b00_00010001110;
storage[820] = 14'b00_00111100110;
storage[821] = -14'b00_00100010111;
storage[822] = -14'b00_01010100001;
storage[823] = -14'b00_00111011010;
storage[824] = -14'b00_00011000010;
storage[825] = 14'b00_00000101000;
storage[826] = 14'b00_00011001011;
storage[827] = -14'b00_00110101001;
storage[828] = -14'b00_00101100010;
storage[829] = 14'b00_00011100001;
storage[830] = -14'b00_01010001010;
storage[831] = -14'b00_00011100000;
storage[832] = -14'b00_00111001000;
storage[833] = -14'b00_01000001011;
storage[834] = 14'b00_00110001000;
storage[835] = 14'b00_10000011010;
storage[836] = -14'b00_00100001000;
storage[837] = 14'b00_01010001111;
storage[838] = -14'b00_00100000000;
storage[839] = -14'b00_01001100000;
storage[840] = 14'b10_00100010000;
storage[841] = -14'b00_00110000100;
storage[842] = -14'b00_01011011010;
storage[843] = -14'b00_01011110010;
storage[844] = -14'b00_01100111001;
storage[845] = -14'b00_00110000111;
storage[846] = 14'b00_00111001010;
storage[847] = -14'b00_10111010010;
storage[848] = -14'b00_00111001100;
storage[849] = 14'b00_00101101101;
storage[850] = -14'b00_00111100010;
storage[851] = -14'b00_00011100000;
storage[852] = 14'b00_00000110110;
storage[853] = 14'b00_00100011010;
storage[854] = 14'b00_00000101111;
storage[855] = 14'b00_00010101010;
storage[856] = 14'b00_00100101000;
storage[857] = 14'b00_01111011000;
storage[858] = 14'b00_00000100000;
storage[859] = -14'b00_01101110011;
storage[860] = -14'b00_00110010000;
storage[861] = 14'b00_01010001100;
storage[862] = -14'b00_00010111100;
storage[863] = -14'b00_00101101111;
storage[864] = 14'b00_01111001100;
storage[865] = 14'b00_00001001101;
storage[866] = -14'b00_01100001000;
storage[867] = 14'b00_00001110011;
storage[868] = -14'b00_00011010011;
storage[869] = -14'b00_01101010001;
storage[870] = 14'b00_00001001011;
storage[871] = 14'b00_00010001111;
storage[872] = 14'b00_00101110000;
storage[873] = 14'b00_00111111000;
storage[874] = -14'b00_01010110011;
storage[875] = -14'b00_00010100111;
storage[876] = 14'b00_01100001100;
storage[877] = 14'b00_01011111000;
storage[878] = -14'b00_01010111100;
storage[879] = 14'b00_00100100111;
storage[880] = -14'b00_00001011100;
storage[881] = -14'b00_10011110101;
storage[882] = 14'b00_10000101010;
storage[883] = -14'b00_00101100011;
storage[884] = -14'b00_01001010100;
storage[885] = -14'b00_00000110011;
storage[886] = -14'b00_01100000110;
storage[887] = 14'b00_00010101101;
//conv4.depthwise.depthwise.weight
storage[888] = -14'b00_01101010100;
storage[889] = -14'b00_00110001100;
storage[890] = -14'b00_01011011001;
storage[891] = 14'b00_00010100010;
storage[892] = -14'b00_00110000101;
storage[893] = -14'b00_01011010111;
storage[894] = -14'b00_01010000110;
storage[895] = 14'b00_00100101000;
storage[896] = -14'b00_01111101001;
storage[897] = 14'b00_00101101111;
storage[898] = 14'b00_00011011111;
storage[899] = 14'b00_01110010001;
storage[900] = 14'b00_00111010101;
storage[901] = -14'b00_00101101001;
storage[902] = 14'b00_01110101101;
storage[903] = 14'b00_00110101000;
storage[904] = 14'b00_00011110001;
storage[905] = 14'b00_00010011101;
storage[906] = 14'b00_00111011011;
storage[907] = -14'b00_00111010110;
storage[908] = 14'b00_00111011000;
storage[909] = -14'b00_00100011010;
storage[910] = -14'b00_00101100100;
storage[911] = -14'b00_00110111010;
storage[912] = -14'b00_00100001110;
storage[913] = -14'b00_01011100010;
storage[914] = -14'b00_00000010000;
storage[915] = -14'b00_01010110110;
storage[916] = 14'b00_00100001011;
storage[917] = 14'b00_00101100110;
storage[918] = -14'b00_00101100011;
storage[919] = -14'b00_00110111101;
storage[920] = -14'b00_01010110111;
storage[921] = -14'b00_00001011011;
storage[922] = 14'b00_00011110010;
storage[923] = 14'b00_00001000000;
storage[924] = -14'b00_00101101111;
storage[925] = -14'b00_00011011110;
storage[926] = 14'b00_01000110100;
storage[927] = 14'b00_00000111011;
storage[928] = -14'b00_00001011110;
storage[929] = 14'b00_00111001001;
storage[930] = 14'b00_00101101110;
storage[931] = 14'b00_01001000011;
storage[932] = 14'b00_00010111101;
storage[933] = -14'b00_01011110000;
storage[934] = -14'b00_00001000000;
storage[935] = 14'b00_01110010100;
storage[936] = -14'b00_01000110100;
storage[937] = 14'b00_01111011110;
storage[938] = 14'b00_01010101011;
storage[939] = -14'b00_00101000010;
storage[940] = 14'b00_01110000011;
storage[941] = 14'b00_01001100100;
//conv4.pointwise.pointwise.weight
storage[942] = 14'b00_01010101111;
storage[943] = 14'b00_00111001111;
storage[944] = -14'b00_10001010010;
storage[945] = -14'b00_00010001110;
storage[946] = 14'b00_00011001000;
storage[947] = 14'b00_00100000001;
storage[948] = -14'b00_00111100101;
storage[949] = 14'b00_00100010101;
storage[950] = 14'b00_00110000011;
storage[951] = 14'b00_01011111111;
storage[952] = -14'b00_01010000000;
storage[953] = 14'b00_00110101000;
storage[954] = 14'b00_01110100101;
storage[955] = 14'b00_01010100101;
storage[956] = -14'b00_10001101001;
storage[957] = -14'b00_01001000110;
storage[958] = 14'b00_00111110110;
storage[959] = 14'b00_10110000110;
//conv5.depthwise.depthwise.weight
storage[960] = -14'b00_01000111011;
storage[961] = -14'b00_01011011000;
storage[962] = 14'b00_00111101010;
storage[963] = -14'b00_01110001010;
storage[964] = -14'b00_01101010000;
storage[965] = -14'b00_00110101010;
storage[966] = -14'b00_00111111001;
storage[967] = -14'b00_01110111100;
storage[968] = -14'b00_00001110000;
storage[969] = 14'b00_10011001001;
storage[970] = 14'b00_01001001110;
storage[971] = 14'b00_00110010000;
storage[972] = -14'b00_01011110011;
storage[973] = -14'b00_01000000100;
storage[974] = -14'b00_00110010010;
storage[975] = -14'b00_00010001000;
storage[976] = 14'b00_00101010010;
storage[977] = 14'b00_00010110001;
storage[978] = 14'b00_00111100110;
storage[979] = -14'b00_01010000101;
storage[980] = 14'b00_00001011101;
storage[981] = -14'b00_00101010000;
storage[982] = -14'b00_01010100101;
storage[983] = 14'b00_00101001101;
storage[984] = -14'b00_01001111110;
storage[985] = -14'b00_01011101111;
storage[986] = 14'b00_00011101000;
//conv5.pointwise.pointwise.weight
storage[987] = -14'b00_00111100001;
storage[988] = 14'b00_10110101000;
storage[989] = -14'b00_01010010001;
	end

	always @(posedge clk) begin
		if(re==1) begin
			datata <= storage[address];
		end
    end
endmodule
